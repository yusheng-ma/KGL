/****************************************************************************
 *                                                                          *
 *  VERILOG VERSION of ORIGINAL NETLIST for c7552                           *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *                                                                          *
 *                Sep 16, 1998                                              *
 *                                                                          *
****************************************************************************/

module c7552g (
        L213, L214, L215, L216, L209, L153, L154, 
        L155, L156, L157, L158, L159, L160, L151, L219, 
        L220, L221, L222, L223, L224, L225, L226, L217, 
        L231, L232, L233, L234, L235, L236, L237, L238, 
        L135, L144, L138, L147, L66, L50, L32, L35, 
        L47, L121, L94, L97, L118, L100, L124, L127, 
        L130, L103, L23, L26, L29, L41, L1486, L1480, 
        L106, L1469, L1462, L2256, L2253, L2247, L2239, L2236, 
        L2230, L2224, L2218, L2211, L4437, L4432, L4427, L4420, 
        L4415, L4410, L4405, L4400, L4394, L3749, L3743, L3737, 
        L3729, L3723, L3717, L3711, L3705, L88, L112, L87, 
        L111, L113, L110, L109, L86, L63, L64, L85, 
        L84, L83, L65, L62, L61, L60, L79, L80, 
        L81, L59, L78, L77, L56, L55, L54, L53, 
        L73, L75, L76, L74, L166, L167, L168, L169, 
        L173, L174, L175, L176, L177, L178, L179, L180, 
        L171, L189, L190, L191, L192, L193, L194, L195, 
        L196, L187, L200, L201, L202, L203, L204, L205, 
        L206, L207, L18, L12, L9, L4526, L89, L38, 
        L4528, L211, L212, L161, L227, L239, L229, L141, 
        L115, L44, L1459, L1496, L1492, L2208, L4393, L3701, 
        L3698, L114, L2204, L1455, L82, L58, L70, L69, 
        L170, L164, L165, L181, L197, L208, L198, L199, 
        L188, L172, L162, L186, L185, L182, L183, L230, 
        L218, L152, L210, L240, L228, L184, L150, L1, 
        L163, L15, L1197, L134, L133, L5, L57, L339,
        L469, L471, L327, L330, L333, L336, L324, 
        L298, L301, L304, L307, L310, L313, L316, L319, 
        L295, L347, L350, L353, L356, L359, L362, L365, 
        L368, L344, L376, L379, L382, L385, L388, L391, 
        L394, L397, L373, L419, L422, L270, L246, L273, 
        L276, L258, L264, L249, L252, L338, L321, L370, 
        L399, L416, L414, L412, L418, L410, L408, L406, 
        L404, L440, L438, L442, L444, L446, L448, L436, 
        L480, L482, L484, L486, L488, L490, L492, L494, 
        L478, L524, L526, L528, L530, L532, L534, L536, 
        L538, L522, L544, L546, L548, L550, L552, L554, 
        L556, L558, L542, L450, L496, L540, L560, L402, 
        L289, L292, L279, L278, L2, L3, L432, L453, 
        L286, L341, L281, L284, L339o);
 
   input
        L213, L214, L215, L216, L209, L153, L154, 
        L155, L156, L157, L158, L159, L160, L151, L219, 
        L220, L221, L222, L223, L224, L225, L226, L217, 
        L231, L232, L233, L234, L235, L236, L237, L238, 
        L135, L144, L138, L147, L66, L50, L32, L35, 
        L47, L121, L94, L97, L118, L100, L124, L127, 
        L130, L103, L23, L26, L29, L41, L1486, L1480, 
        L106, L1469, L1462, L2256, L2253, L2247, L2239, L2236, 
        L2230, L2224, L2218, L2211, L4437, L4432, L4427, L4420, 
        L4415, L4410, L4405, L4400, L4394, L3749, L3743, L3737, 
        L3729, L3723, L3717, L3711, L3705, L88, L112, L87, 
        L111, L113, L110, L109, L86, L63, L64, L85, 
        L84, L83, L65, L62, L61, L60, L79, L80, 
        L81, L59, L78, L77, L56, L55, L54, L53, 
        L73, L75, L76, L74, L166, L167, L168, L169, 
        L173, L174, L175, L176, L177, L178, L179, L180, 
        L171, L189, L190, L191, L192, L193, L194, L195, 
        L196, L187, L200, L201, L202, L203, L204, L205, 
        L206, L207, L18, L12, L9, L4526, L89, L38, 
        L4528, L211, L212, L161, L227, L239, L229, L141, 
        L115, L44, L1459, L1496, L1492, L2208, L4393, L3701, 
        L3698, L114, L2204, L1455, L82, L58, L70, L69, 
        L170, L164, L165, L181, L197, L208, L198, L199, 
        L188, L172, L162, L186, L185, L182, L183, L230, 
        L218, L152, L210, L240, L228, L184, L150, L1, 
        L163, L15, L1197, L134, L133, L5, L57, L339;
 
   output
        L469, L471, L327, L330, L333, L336, L324, 
        L298, L301, L304, L307, L310, L313, L316, L319, 
        L295, L347, L350, L353, L356, L359, L362, L365, 
        L368, L344, L376, L379, L382, L385, L388, L391, 
        L394, L397, L373, L419, L422, L270, L246, L273, 
        L276, L258, L264, L249, L252, L338, L321, L370, 
        L399, L416, L414, L412, L418, L410, L408, L406, 
        L404, L440, L438, L442, L444, L446, L448, L436, 
        L480, L482, L484, L486, L488, L490, L492, L494, 
        L478, L524, L526, L528, L530, L532, L534, L536, 
        L538, L522, L544, L546, L548, L550, L552, L554, 
        L556, L558, L542, L450, L496, L540, L560, L402, 
        L289, L292, L279, L278, L2, L3, L432, L453, 
        L286, L341, L281, L284, L339o;


   assign L339o = L339; 


   buffer U2 ( L1, L2 ); 
   buffer U3 ( L1, L3 ); 
   inv U4 ( L57, L400 ); 
   and2 U5 ( L134, L133, L1184 ); 
   buffer U6 ( L1459, L450 ); 
   buffer U7 ( L1469, L448 ); 
   buffer U8 ( L1480, L444 ); 
   buffer U9 ( L1486, L442 ); 
   buffer U10 ( L1492, L440 ); 
   buffer U11 ( L1496, L438 ); 
   and4 U12 ( L162, L172, L188, L199, L1501 ); 
   buffer U13 ( L2208, L496 ); 
   buffer U14 ( L2218, L494 ); 
   buffer U15 ( L2224, L492 ); 
   buffer U16 ( L2230, L490 ); 
   buffer U17 ( L2236, L488 ); 
   buffer U18 ( L2239, L486 ); 
   buffer U19 ( L2247, L484 ); 
   buffer U20 ( L2253, L482 ); 
   buffer U21 ( L2256, L480 ); 
   and4 U22 ( L150, L184, L228, L240, L2857 ); 
   buffer U23 ( L3698, L560 ); 
   buffer U24 ( L3701, L542 ); 
   buffer U25 ( L3705, L558 ); 
   buffer U26 ( L3711, L556 ); 
   buffer U27 ( L3717, L554 ); 
   buffer U28 ( L3723, L552 ); 
   buffer U29 ( L3729, L550 ); 
   buffer U30 ( L3737, L548 ); 
   buffer U31 ( L3743, L546 ); 
   buffer U32 ( L3749, L544 ); 
   buffer U33 ( L4393, L540 ); 
   buffer U34 ( L4400, L538 ); 
   buffer U35 ( L4405, L536 ); 
   buffer U36 ( L4410, L534 ); 
   buffer U37 ( L4415, L532 ); 
   buffer U38 ( L4420, L530 ); 
   buffer U39 ( L4427, L528 ); 
   buffer U40 ( L4432, L526 ); 
   buffer U41 ( L4437, L524 ); 
   and4 U42 ( L183, L182, L185, L186, L4442 ); 
   and4 U43 ( L210, L152, L218, L230, L4514 ); 
   inv U44 ( L15, L279 ); 
   inv U45 ( L5, L401 ); 
   buffer U46 ( L1, L573 ); 
   inv U47 ( L5, L574 ); 
   inv U48 ( L5, L575 ); 
   inv U49 ( L2236, L1178 ); 
   inv U50 ( L2253, L1186 ); 
   inv U51 ( L2256, L1192 ); 
   buffer U52 ( L38, L1198 ); 
   buffer U53 ( L15, L1205 ); 
   nand2 U54 ( L12, L9, L1206 ); 
   nand2 U55 ( L12, L9, L1207 ); 
   buffer U56 ( L38, L1210 ); 
   inv U57 ( L1455, L1458 ); 
   inv U58 ( L1459, L1461 ); 
   buffer U59 ( L1462, L436 ); 
   inv U60 ( L1462, L1464 ); 
   inv U61 ( L1469, L1471 ); 
   buffer U62 ( L106, L1475 ); 
   inv U63 ( L1480, L1482 ); 
   inv U64 ( L1486, L1488 ); 
   inv U65 ( L1492, L1495 ); 
   inv U66 ( L1496, L1499 ); 
   inv U67 ( L106, L1500 ); 
   buffer U68 ( L18, L1503 ); 
   buffer U69 ( L18, L1512 ); 
   and2 U70 ( L4528, L1492, L1518 ); 
   buffer U71 ( L18, L1524 ); 
   inv U72 ( L18, L1535 ); 
   nand2 U73 ( L4528, L1496, L1541 ); 
   inv U74 ( L2204, L2207 ); 
   inv U75 ( L2208, L2210 ); 
   buffer U76 ( L2211, L478 ); 
   inv U77 ( L2211, L2213 ); 
   inv U78 ( L2218, L2220 ); 
   inv U79 ( L2224, L2226 ); 
   inv U80 ( L2230, L2232 ); 
   inv U81 ( L2236, L2238 ); 
   inv U82 ( L2239, L2241 ); 
   inv U83 ( L2247, L2249 ); 
   inv U84 ( L2253, L2255 ); 
   inv U85 ( L2256, L2258 ); 
   buffer U86 ( L4526, L2828 ); 
   inv U87 ( L3698, L3700 ); 
   inv U88 ( L3701, L3703 ); 
   inv U89 ( L3705, L3707 ); 
   inv U90 ( L3711, L3713 ); 
   inv U91 ( L3717, L3719 ); 
   inv U92 ( L3723, L3725 ); 
   inv U93 ( L3729, L3731 ); 
   inv U94 ( L3737, L3739 ); 
   inv U95 ( L3743, L3745 ); 
   inv U96 ( L3749, L3751 ); 
   inv U97 ( L4393, L4121 ); 
   buffer U98 ( L4394, L522 ); 
   inv U99 ( L4394, L4396 ); 
   inv U100 ( L4400, L4402 ); 
   inv U101 ( L4405, L4407 ); 
   inv U102 ( L4410, L4412 ); 
   inv U103 ( L4415, L4417 ); 
   inv U104 ( L4420, L4422 ); 
   inv U105 ( L4427, L4429 ); 
   inv U106 ( L4432, L4434 ); 
   inv U107 ( L4437, L4439 ); 
   buffer U108 ( L4526, L4833 ); 
   nand2 U109 ( L400, L401, L402 ); 
   inv U110 ( L2857, L404 ); 
   inv U111 ( L4514, L406 ); 
   inv U112 ( L4442, L408 ); 
   inv U113 ( L1501, L410 ); 
   and2 U114 ( L2857, L4514, L2876 ); 
   and2 U115 ( L4442, L1501, L2878 ); 
   buffer U116 ( L573, L432 ); 
   buffer U117 ( L1475, L446 ); 
   inv U118 ( L1518, L1519 ); 
   and2 U119 ( L4528, L1458, L2871 ); 
   nand2 U120 ( L4528, L2207, L2883 ); 
   and2 U121 ( L1184, L575, L280 ); 
   nand2 U122 ( L1197, L574, L284 ); 
   inv U123 ( L1205, L286 ); 
   nand2 U124 ( L1197, L574, L289 ); 
   nand2 U125 ( L1184, L575, L292 ); 
   inv U126 ( L1205, L341 ); 
   inv U127 ( L4833, L4839 ); 
   buffer U128 ( L573, L572 ); 
   buffer U129 ( L1206, L581 ); 
   buffer U130 ( L1512, L587 ); 
   buffer U131 ( L1206, L601 ); 
   buffer U132 ( L1512, L606 ); 
   buffer U133 ( L1206, L650 ); 
   buffer U134 ( L1512, L657 ); 
   buffer U135 ( L1207, L671 ); 
   buffer U136 ( L1503, L678 ); 
   and2 U137 ( L1541, L1198, L777 ); 
   and2 U138 ( L1541, L1198, L1115 ); 
   buffer U139 ( L1512, L1336 ); 
   buffer U140 ( L1503, L1350 ); 
   inv U141 ( L1475, L1477 ); 
   inv U142 ( L1503, L1507 ); 
   inv U143 ( L1512, L1514 ); 
   inv U144 ( L1524, L1530 ); 
   buffer U145 ( L1535, L2259 ); 
   inv U146 ( L2828, L2833 ); 
   inv U147 ( L2871, L2872 ); 
   buffer U148 ( L1207, L2886 ); 
   buffer U149 ( L1503, L2892 ); 
   buffer U150 ( L1207, L2905 ); 
   buffer U151 ( L1503, L2909 ); 
   buffer U152 ( L1524, L3622 ); 
   buffer U153 ( L1524, L3635 ); 
   buffer U154 ( L1535, L3755 ); 
   buffer U155 ( L1524, L4640 ); 
   buffer U156 ( L1524, L4653 ); 
   buffer U157 ( L1541, L4873 ); 
   buffer U158 ( L1198, L4876 ); 
   buffer U159 ( L1488, L4881 ); 
   buffer U160 ( L1482, L4889 ); 
   buffer U161 ( L1471, L4905 ); 
   buffer U162 ( L1198, L4916 ); 
   buffer U163 ( L1464, L4921 ); 
   buffer U164 ( L1541, L5175 ); 
   buffer U165 ( L1198, L5178 ); 
   buffer U166 ( L1198, L5186 ); 
   buffer U167 ( L1488, L5191 ); 
   buffer U168 ( L1482, L5199 ); 
   buffer U169 ( L1471, L5215 ); 
   buffer U170 ( L1464, L5223 ); 
   buffer U171 ( L1192, L5393 ); 
   buffer U172 ( L1186, L5401 ); 
   buffer U173 ( L2249, L5409 ); 
   buffer U174 ( L1178, L5417 ); 
   buffer U175 ( L2232, L5425 ); 
   buffer U176 ( L2226, L5433 ); 
   buffer U177 ( L2220, L5441 ); 
   buffer U178 ( L2241, L5449 ); 
   buffer U179 ( L2213, L5457 ); 
   buffer U180 ( L1192, L5745 ); 
   buffer U181 ( L1186, L5753 ); 
   buffer U182 ( L2249, L5761 ); 
   buffer U183 ( L2241, L5769 ); 
   buffer U184 ( L1178, L5777 ); 
   buffer U185 ( L2232, L5785 ); 
   buffer U186 ( L2226, L5793 ); 
   buffer U187 ( L2220, L5801 ); 
   buffer U188 ( L2213, L5809 ); 
   buffer U189 ( L3751, L5865 ); 
   buffer U190 ( L3745, L5873 ); 
   buffer U191 ( L3739, L5881 ); 
   buffer U192 ( L3731, L5889 ); 
   buffer U193 ( L3725, L5897 ); 
   buffer U194 ( L3719, L5905 ); 
   buffer U195 ( L3713, L5913 ); 
   buffer U196 ( L3707, L5921 ); 
   buffer U197 ( L3751, L5985 ); 
   buffer U198 ( L3745, L5993 ); 
   buffer U199 ( L3739, L6001 ); 
   buffer U200 ( L3725, L6009 ); 
   buffer U201 ( L3719, L6017 ); 
   buffer U202 ( L3713, L6025 ); 
   buffer U203 ( L3707, L6033 ); 
   buffer U204 ( L3731, L6041 ); 
   buffer U205 ( L1210, L6514 ); 
   buffer U206 ( L1210, L6554 ); 
   buffer U207 ( L4439, L6567 ); 
   buffer U208 ( L4434, L6575 ); 
   buffer U209 ( L4429, L6583 ); 
   buffer U210 ( L4422, L6591 ); 
   buffer U211 ( L4417, L6599 ); 
   buffer U212 ( L4412, L6607 ); 
   buffer U213 ( L4407, L6615 ); 
   buffer U214 ( L4402, L6623 ); 
   buffer U215 ( L4396, L6631 ); 
   buffer U216 ( L4439, L6853 ); 
   buffer U217 ( L4434, L6861 ); 
   buffer U218 ( L4429, L6869 ); 
   buffer U219 ( L4417, L6877 ); 
   buffer U220 ( L4412, L6885 ); 
   buffer U221 ( L4407, L6893 ); 
   buffer U222 ( L4402, L6901 ); 
   buffer U223 ( L4422, L6909 ); 
   buffer U224 ( L4396, L6917 ); 
   inv U225 ( L280, L281 ); 
   buffer U226 ( L572, L453 ); 
   and2 U227 ( L1519, L1198, L784 ); 
   and2 U228 ( L1198, L1519, L1014 ); 
   and2 U229 ( L2883, L1210, L3221 ); 
   buffer U230 ( L1519, L4913 ); 
   nor2 U231 ( L1519, L1198, L4929 ); 
   buffer U232 ( L1519, L5183 ); 
   nor2 U233 ( L1198, L1519, L5231 ); 
   buffer U234 ( L2883, L6511 ); 
   and2 U235 ( L163, L572, L278 ); 
   and2 U236 ( L170, L587, L615 ); 
   inv U237 ( L587, L594 ); 
   inv U238 ( L606, L611 ); 
   and2 U239 ( L169, L587, L617 ); 
   and2 U240 ( L168, L587, L619 ); 
   and2 U241 ( L167, L587, L621 ); 
   and2 U242 ( L166, L606, L623 ); 
   and2 U243 ( L165, L606, L625 ); 
   and2 U244 ( L164, L606, L627 ); 
   inv U245 ( L657, L664 ); 
   inv U246 ( L678, L685 ); 
   and2 U247 ( L177, L657, L691 ); 
   and2 U248 ( L176, L657, L693 ); 
   and2 U249 ( L175, L657, L695 ); 
   and2 U250 ( L174, L657, L697 ); 
   and2 U251 ( L173, L657, L699 ); 
   and2 U252 ( L157, L678, L701 ); 
   and2 U253 ( L156, L678, L703 ); 
   and2 U254 ( L155, L678, L705 ); 
   and2 U255 ( L154, L678, L707 ); 
   and2 U256 ( L153, L678, L709 ); 
   inv U257 ( L4873, L4879 ); 
   inv U258 ( L4876, L4880 ); 
   inv U259 ( L4881, L4887 ); 
   inv U260 ( L4889, L4895 ); 
   inv U261 ( L4905, L4911 ); 
   inv U262 ( L4916, L4920 ); 
   inv U263 ( L4921, L4927 ); 
   inv U264 ( L5175, L5181 ); 
   inv U265 ( L5178, L5182 ); 
   inv U266 ( L5186, L5190 ); 
   inv U267 ( L5191, L5197 ); 
   inv U268 ( L5199, L5205 ); 
   inv U269 ( L5215, L5221 ); 
   inv U270 ( L5223, L5229 ); 
   inv U271 ( L1336, L1343 ); 
   inv U272 ( L1350, L1357 ); 
   and2 U273 ( L181, L1336, L1364 ); 
   and2 U274 ( L171, L1336, L1366 ); 
   and2 U275 ( L180, L1336, L1368 ); 
   and2 U276 ( L179, L1336, L1370 ); 
   and2 U277 ( L178, L1336, L1372 ); 
   and2 U278 ( L161, L1350, L1374 ); 
   and2 U279 ( L151, L1350, L1376 ); 
   and2 U280 ( L160, L1350, L1378 ); 
   and2 U281 ( L159, L1350, L1380 ); 
   and2 U282 ( L158, L1350, L1382 ); 
   inv U283 ( L5393, L5399 ); 
   inv U284 ( L5401, L5407 ); 
   inv U285 ( L5409, L5415 ); 
   inv U286 ( L5417, L5423 ); 
   inv U287 ( L5425, L5431 ); 
   inv U288 ( L5433, L5439 ); 
   inv U289 ( L5441, L5447 ); 
   inv U290 ( L5449, L5455 ); 
   inv U291 ( L5457, L5463 ); 
   inv U292 ( L5745, L5751 ); 
   inv U293 ( L5753, L5759 ); 
   inv U294 ( L5761, L5767 ); 
   inv U295 ( L5769, L5775 ); 
   inv U296 ( L5777, L5783 ); 
   inv U297 ( L5785, L5791 ); 
   inv U298 ( L5793, L5799 ); 
   inv U299 ( L5801, L5807 ); 
   inv U300 ( L5809, L5815 ); 
   buffer U301 ( L1514, L2019 ); 
   buffer U302 ( L1507, L2032 ); 
   buffer U303 ( L1514, L2117 ); 
   buffer U304 ( L1507, L2130 ); 
   inv U305 ( L2259, L2266 ); 
   buffer U306 ( L1507, L2272 ); 
   and2 U307 ( L44, L2259, L2286 ); 
   and2 U308 ( L41, L2259, L2288 ); 
   and2 U309 ( L29, L2259, L2290 ); 
   and2 U310 ( L26, L2259, L2292 ); 
   and2 U311 ( L23, L2259, L2294 ); 
   inv U312 ( L5865, L5871 ); 
   inv U313 ( L5873, L5879 ); 
   inv U314 ( L5881, L5887 ); 
   inv U315 ( L5889, L5895 ); 
   inv U316 ( L5897, L5903 ); 
   inv U317 ( L5905, L5911 ); 
   inv U318 ( L5913, L5919 ); 
   inv U319 ( L5921, L5927 ); 
   inv U320 ( L5985, L5991 ); 
   inv U321 ( L5993, L5999 ); 
   inv U322 ( L6001, L6007 ); 
   inv U323 ( L6009, L6015 ); 
   inv U324 ( L6017, L6023 ); 
   inv U325 ( L6025, L6031 ); 
   inv U326 ( L6033, L6039 ); 
   inv U327 ( L6041, L6047 ); 
   inv U328 ( L2892, L2899 ); 
   inv U329 ( L2909, L2914 ); 
   and2 U330 ( L209, L2892, L2919 ); 
   and2 U331 ( L216, L2892, L2921 ); 
   and2 U332 ( L215, L2892, L2923 ); 
   and2 U333 ( L214, L2892, L2925 ); 
   and2 U334 ( L213, L2909, L2927 ); 
   and2 U335 ( L212, L2909, L2929 ); 
   and2 U336 ( L211, L2909, L2931 ); 
   inv U337 ( L6514, L6518 ); 
   and2 U338 ( L2872, L1210, L3173 ); 
   inv U339 ( L6554, L6558 ); 
   inv U340 ( L6567, L6573 ); 
   inv U341 ( L6575, L6581 ); 
   inv U342 ( L6583, L6589 ); 
   inv U343 ( L6591, L6597 ); 
   inv U344 ( L6599, L6605 ); 
   inv U345 ( L6607, L6613 ); 
   inv U346 ( L6615, L6621 ); 
   inv U347 ( L6623, L6629 ); 
   inv U348 ( L6631, L6637 ); 
   inv U349 ( L3622, L3629 ); 
   inv U350 ( L3635, L3642 ); 
   and2 U351 ( L1461, L3622, L3649 ); 
   and2 U352 ( L1464, L3622, L3651 ); 
   and2 U353 ( L1471, L3622, L3653 ); 
   and2 U354 ( L1500, L3622, L3655 ); 
   and2 U355 ( L1482, L3622, L3657 ); 
   and2 U356 ( L1488, L3635, L3659 ); 
   and2 U357 ( L1495, L3635, L3661 ); 
   and2 U358 ( L1499, L3635, L3663 ); 
   inv U359 ( L3755, L3762 ); 
   buffer U360 ( L1507, L3768 ); 
   and2 U361 ( L47, L3755, L3782 ); 
   and2 U362 ( L35, L3755, L3784 ); 
   and2 U363 ( L32, L3755, L3786 ); 
   and2 U364 ( L50, L3755, L3788 ); 
   and2 U365 ( L66, L3755, L3790 ); 
   inv U366 ( L6853, L6859 ); 
   inv U367 ( L6861, L6867 ); 
   inv U368 ( L6869, L6875 ); 
   inv U369 ( L6877, L6883 ); 
   inv U370 ( L6885, L6891 ); 
   inv U371 ( L6893, L6899 ); 
   inv U372 ( L6901, L6907 ); 
   inv U373 ( L6909, L6915 ); 
   inv U374 ( L6917, L6923 ); 
   buffer U375 ( L1530, L4094 ); 
   buffer U376 ( L1530, L4107 ); 
   buffer U377 ( L1530, L4444 ); 
   buffer U378 ( L1530, L4457 ); 
   inv U379 ( L4640, L4647 ); 
   inv U380 ( L4653, L4660 ); 
   and2 U381 ( L2210, L4640, L4667 ); 
   and2 U382 ( L2213, L4640, L4669 ); 
   and2 U383 ( L2220, L4640, L4671 ); 
   and2 U384 ( L2226, L4640, L4673 ); 
   and2 U385 ( L2232, L4640, L4675 ); 
   and2 U386 ( L2238, L4653, L4677 ); 
   and2 U387 ( L2241, L4653, L4679 ); 
   and2 U388 ( L2249, L4653, L4681 ); 
   and2 U389 ( L2255, L4653, L4683 ); 
   and2 U390 ( L2258, L4653, L4685 ); 
   buffer U391 ( L1477, L4897 ); 
   buffer U392 ( L1477, L5207 ); 
   buffer U393 ( L2872, L6551 ); 
   nand2 U394 ( L4876, L4879, L763 ); 
   nand2 U395 ( L4873, L4880, L764 ); 
   inv U396 ( L4913, L4919 ); 
   nand2 U397 ( L4913, L4920, L886 ); 
   nand2 U398 ( L5178, L5181, L1005 ); 
   nand2 U399 ( L5175, L5182, L1006 ); 
   inv U400 ( L5183, L5189 ); 
   nand2 U401 ( L5183, L5190, L1018 ); 
   inv U402 ( L5231, L5237 ); 
   inv U403 ( L6511, L6517 ); 
   nand2 U404 ( L6511, L6518, L3169 ); 
   inv U405 ( L4929, L4935 ); 
   buffer U406 ( L784, L4970 ); 
   buffer U407 ( L1014, L5239 ); 
   or2 U408 ( L594, L615, L577 ); 
   or2 U409 ( L594, L587, L616 ); 
   or2 U410 ( L594, L617, L618 ); 
   or2 U411 ( L594, L619, L620 ); 
   or2 U412 ( L594, L621, L622 ); 
   or2 U413 ( L611, L623, L624 ); 
   or2 U414 ( L611, L625, L626 ); 
   or2 U415 ( L611, L627, L628 ); 
   or2 U416 ( L664, L691, L692 ); 
   or2 U417 ( L664, L693, L694 ); 
   or2 U418 ( L664, L695, L696 ); 
   or2 U419 ( L664, L697, L698 ); 
   or2 U420 ( L664, L699, L700 ); 
   or2 U421 ( L685, L701, L702 ); 
   or2 U422 ( L685, L703, L704 ); 
   or2 U423 ( L685, L705, L706 ); 
   or2 U424 ( L685, L707, L708 ); 
   or2 U425 ( L685, L709, L710 ); 
   nand2 U426 ( L763, L764, L765 ); 
   inv U427 ( L4897, L4903 ); 
   nand2 U428 ( L4916, L4919, L885 ); 
   nand2 U429 ( L1005, L1006, L1007 ); 
   nand2 U430 ( L5186, L5189, L1017 ); 
   inv U431 ( L5207, L5213 ); 
   and2 U432 ( L141, L1343, L1363 ); 
   and2 U433 ( L147, L1343, L1365 ); 
   and2 U434 ( L138, L1343, L1367 ); 
   and2 U435 ( L144, L1343, L1369 ); 
   and2 U436 ( L135, L1343, L1371 ); 
   and2 U437 ( L141, L1357, L1373 ); 
   and2 U438 ( L147, L1357, L1375 ); 
   and2 U439 ( L138, L1357, L1377 ); 
   and2 U440 ( L144, L1357, L1379 ); 
   and2 U441 ( L135, L1357, L1381 ); 
   inv U442 ( L2019, L2026 ); 
   inv U443 ( L2032, L2039 ); 
   and2 U444 ( L103, L2019, L2046 ); 
   and2 U445 ( L130, L2019, L2048 ); 
   and2 U446 ( L127, L2019, L2050 ); 
   and2 U447 ( L124, L2019, L2052 ); 
   and2 U448 ( L100, L2019, L2054 ); 
   and2 U449 ( L103, L2032, L2056 ); 
   and2 U450 ( L130, L2032, L2058 ); 
   and2 U451 ( L127, L2032, L2060 ); 
   and2 U452 ( L124, L2032, L2062 ); 
   and2 U453 ( L100, L2032, L2064 ); 
   inv U454 ( L2117, L2124 ); 
   inv U455 ( L2130, L2137 ); 
   and2 U456 ( L115, L2117, L2144 ); 
   and2 U457 ( L118, L2117, L2146 ); 
   and2 U458 ( L97, L2117, L2148 ); 
   and2 U459 ( L94, L2117, L2150 ); 
   and2 U460 ( L121, L2117, L2152 ); 
   and2 U461 ( L115, L2130, L2154 ); 
   and2 U462 ( L118, L2130, L2156 ); 
   and2 U463 ( L97, L2130, L2158 ); 
   and2 U464 ( L94, L2130, L2160 ); 
   and2 U465 ( L121, L2130, L2162 ); 
   inv U466 ( L2272, L2279 ); 
   and2 U467 ( L208, L2266, L2285 ); 
   and2 U468 ( L198, L2266, L2287 ); 
   and2 U469 ( L207, L2266, L2289 ); 
   and2 U470 ( L206, L2266, L2291 ); 
   and2 U471 ( L205, L2266, L2293 ); 
   and2 U472 ( L44, L2272, L2296 ); 
   and2 U473 ( L41, L2272, L2298 ); 
   and2 U474 ( L29, L2272, L2300 ); 
   and2 U475 ( L26, L2272, L2302 ); 
   and2 U476 ( L23, L2272, L2304 ); 
   or2 U477 ( L2899, L2892, L2918 ); 
   or2 U478 ( L2899, L2919, L2920 ); 
   or2 U479 ( L2899, L2921, L2922 ); 
   or2 U480 ( L2899, L2923, L2924 ); 
   or2 U481 ( L2899, L2925, L2926 ); 
   or2 U482 ( L2914, L2927, L2928 ); 
   or2 U483 ( L2914, L2929, L2930 ); 
   or2 U484 ( L2914, L2931, L2932 ); 
   nand2 U485 ( L6514, L6517, L3168 ); 
   inv U486 ( L6551, L6557 ); 
   nand2 U487 ( L6551, L6558, L3211 ); 
   and2 U488 ( L114, L3629, L3648 ); 
   and2 U489 ( L113, L3629, L3650 ); 
   and2 U490 ( L111, L3629, L3652 ); 
   and2 U491 ( L87, L3629, L3654 ); 
   and2 U492 ( L112, L3629, L3656 ); 
   and2 U493 ( L88, L3642, L3658 ); 
   and2 U494 ( L1455, L3642, L3660 ); 
   and2 U495 ( L2204, L3642, L3662 ); 
   and2 U496 ( L3703, L3642, L3665 ); 
   and2 U497 ( L70, L3642, L3666 ); 
   inv U498 ( L3768, L3775 ); 
   and2 U499 ( L193, L3762, L3781 ); 
   and2 U500 ( L192, L3762, L3783 ); 
   and2 U501 ( L191, L3762, L3785 ); 
   and2 U502 ( L190, L3762, L3787 ); 
   and2 U503 ( L189, L3762, L3789 ); 
   and2 U504 ( L47, L3768, L3792 ); 
   and2 U505 ( L35, L3768, L3794 ); 
   and2 U506 ( L32, L3768, L3796 ); 
   and2 U507 ( L50, L3768, L3798 ); 
   and2 U508 ( L66, L3768, L3800 ); 
   inv U509 ( L4094, L4101 ); 
   inv U510 ( L4107, L4114 ); 
   and2 U511 ( L58, L4094, L4123 ); 
   and2 U512 ( L77, L4094, L4126 ); 
   and2 U513 ( L78, L4094, L4129 ); 
   and2 U514 ( L59, L4094, L4132 ); 
   and2 U515 ( L81, L4094, L4135 ); 
   and2 U516 ( L80, L4107, L4138 ); 
   and2 U517 ( L79, L4107, L4141 ); 
   and2 U518 ( L60, L4107, L4144 ); 
   and2 U519 ( L61, L4107, L4147 ); 
   and2 U520 ( L62, L4107, L4150 ); 
   inv U521 ( L4444, L4451 ); 
   inv U522 ( L4457, L4464 ); 
   and2 U523 ( L69, L4444, L4471 ); 
   and2 U524 ( L70, L4444, L4473 ); 
   and2 U525 ( L74, L4444, L4475 ); 
   and2 U526 ( L76, L4444, L4477 ); 
   and2 U527 ( L75, L4444, L4479 ); 
   and2 U528 ( L73, L4457, L4481 ); 
   and2 U529 ( L53, L4457, L4483 ); 
   and2 U530 ( L54, L4457, L4485 ); 
   and2 U531 ( L55, L4457, L4487 ); 
   and2 U532 ( L56, L4457, L4489 ); 
   and2 U533 ( L82, L4647, L4666 ); 
   and2 U534 ( L65, L4647, L4668 ); 
   and2 U535 ( L83, L4647, L4670 ); 
   and2 U536 ( L84, L4647, L4672 ); 
   and2 U537 ( L85, L4647, L4674 ); 
   and2 U538 ( L64, L4660, L4676 ); 
   and2 U539 ( L63, L4660, L4678 ); 
   and2 U540 ( L86, L4660, L4680 ); 
   and2 U541 ( L109, L4660, L4682 ); 
   and2 U542 ( L110, L4660, L4684 ); 
   and2 U543 ( L577, L581, L579 ); 
   and2 U544 ( L616, L581, L629 ); 
   and2 U545 ( L618, L581, L633 ); 
   and2 U546 ( L620, L581, L637 ); 
   and2 U547 ( L622, L581, L641 ); 
   and2 U548 ( L624, L601, L645 ); 
   and2 U549 ( L692, L650, L711 ); 
   and2 U550 ( L694, L650, L715 ); 
   and2 U551 ( L696, L650, L719 ); 
   and2 U552 ( L698, L650, L723 ); 
   and2 U553 ( L700, L650, L727 ); 
   and2 U554 ( L702, L671, L731 ); 
   and2 U555 ( L704, L671, L737 ); 
   and2 U556 ( L706, L671, L745 ); 
   and2 U557 ( L708, L671, L751 ); 
   and2 U558 ( L710, L671, L757 ); 
   nand2 U559 ( L885, L886, L887 ); 
   nand2 U560 ( L1017, L1018, L1019 ); 
   inv U561 ( L5239, L5245 ); 
   or2 U562 ( L1365, L1366, L1383 ); 
   or2 U563 ( L1367, L1368, L1387 ); 
   or2 U564 ( L1369, L1370, L1391 ); 
   or2 U565 ( L1371, L1372, L1395 ); 
   or2 U566 ( L1375, L1376, L1399 ); 
   or2 U567 ( L1377, L1378, L1406 ); 
   or2 U568 ( L1379, L1380, L1412 ); 
   or2 U569 ( L1381, L1382, L1418 ); 
   or2 U570 ( L2287, L2288, L2305 ); 
   or2 U571 ( L2289, L2290, L2308 ); 
   or2 U572 ( L2291, L2292, L2312 ); 
   or2 U573 ( L2293, L2294, L2316 ); 
   and2 U574 ( L2920, L2886, L2933 ); 
   and2 U575 ( L2922, L2886, L2938 ); 
   and2 U576 ( L2924, L2886, L2942 ); 
   and2 U577 ( L2926, L2886, L2946 ); 
   and2 U578 ( L2928, L2905, L2950 ); 
   nand2 U579 ( L3168, L3169, L3170 ); 
   nand2 U580 ( L6554, L6557, L3210 ); 
   or2 U581 ( L3650, L3651, L3667 ); 
   or2 U582 ( L3652, L3653, L3670 ); 
   or2 U583 ( L3654, L3655, L3673 ); 
   or2 U584 ( L3656, L3657, L3676 ); 
   or2 U585 ( L3658, L3659, L3679 ); 
   or2 U586 ( L3665, L3635, L3682 ); 
   or2 U587 ( L3666, L3635, L3686 ); 
   or2 U588 ( L3781, L3782, L3801 ); 
   or2 U589 ( L3783, L3784, L3804 ); 
   or2 U590 ( L3785, L3786, L3807 ); 
   or2 U591 ( L3787, L3788, L3810 ); 
   or2 U592 ( L3789, L3790, L3813 ); 
   and2 U593 ( L2918, L2886, L4525 ); 
   or2 U594 ( L4668, L4669, L4686 ); 
   or2 U595 ( L4670, L4671, L4689 ); 
   or2 U596 ( L4672, L4673, L4692 ); 
   or2 U597 ( L4674, L4675, L4695 ); 
   or2 U598 ( L4676, L4677, L4698 ); 
   or2 U599 ( L4678, L4679, L4701 ); 
   or2 U600 ( L4680, L4681, L4704 ); 
   or2 U601 ( L4682, L4683, L4707 ); 
   or2 U602 ( L4684, L4685, L4710 ); 
   inv U603 ( L4970, L4976 ); 
   and2 U604 ( L2932, L2905, L5271 ); 
   and2 U605 ( L2930, L2905, L5274 ); 
   and2 U606 ( L628, L601, L5305 ); 
   and2 U607 ( L626, L601, L5308 ); 
   or2 U608 ( L1373, L1374, L5318 ); 
   or2 U609 ( L3648, L3649, L6690 ); 
   or2 U610 ( L3662, L3663, L6711 ); 
   or2 U611 ( L3660, L3661, L6714 ); 
   or2 U612 ( L2285, L2286, L7252 ); 
   or2 U613 ( L1363, L1364, L7296 ); 
   or2 U614 ( L4666, L4667, L7466 ); 
   and2 U615 ( L765, L784, L907 ); 
   and2 U616 ( L765, L784, L913 ); 
   and2 U617 ( L765, L784, L915 ); 
   and2 U618 ( L765, L784, L916 ); 
   and2 U619 ( L1007, L1014, L1116 ); 
   and2 U620 ( L204, L2026, L2045 ); 
   and2 U621 ( L203, L2026, L2047 ); 
   and2 U622 ( L202, L2026, L2049 ); 
   and2 U623 ( L201, L2026, L2051 ); 
   and2 U624 ( L200, L2026, L2053 ); 
   and2 U625 ( L235, L2039, L2055 ); 
   and2 U626 ( L234, L2039, L2057 ); 
   and2 U627 ( L233, L2039, L2059 ); 
   and2 U628 ( L232, L2039, L2061 ); 
   and2 U629 ( L231, L2039, L2063 ); 
   and2 U630 ( L197, L2124, L2143 ); 
   and2 U631 ( L187, L2124, L2145 ); 
   and2 U632 ( L196, L2124, L2147 ); 
   and2 U633 ( L195, L2124, L2149 ); 
   and2 U634 ( L194, L2124, L2151 ); 
   and2 U635 ( L227, L2137, L2153 ); 
   and2 U636 ( L217, L2137, L2155 ); 
   and2 U637 ( L226, L2137, L2157 ); 
   and2 U638 ( L225, L2137, L2159 ); 
   and2 U639 ( L224, L2137, L2161 ); 
   and2 U640 ( L239, L2279, L2295 ); 
   and2 U641 ( L229, L2279, L2297 ); 
   and2 U642 ( L238, L2279, L2299 ); 
   and2 U643 ( L237, L2279, L2301 ); 
   and2 U644 ( L236, L2279, L2303 ); 
   nand2 U645 ( L3210, L3211, L3212 ); 
   and2 U646 ( L223, L3775, L3791 ); 
   and2 U647 ( L222, L3775, L3793 ); 
   and2 U648 ( L221, L3775, L3795 ); 
   and2 U649 ( L220, L3775, L3797 ); 
   and2 U650 ( L219, L3775, L3799 ); 
   and2 U651 ( L4121, L4101, L4122 ); 
   and2 U652 ( L4396, L4101, L4125 ); 
   and2 U653 ( L4402, L4101, L4128 ); 
   and2 U654 ( L4407, L4101, L4131 ); 
   and2 U655 ( L4412, L4101, L4134 ); 
   and2 U656 ( L4417, L4114, L4137 ); 
   and2 U657 ( L4422, L4114, L4140 ); 
   and2 U658 ( L4429, L4114, L4143 ); 
   and2 U659 ( L4434, L4114, L4146 ); 
   and2 U660 ( L4439, L4114, L4149 ); 
   and2 U661 ( L3700, L4451, L4470 ); 
   and2 U662 ( L3703, L4451, L4472 ); 
   and2 U663 ( L3707, L4451, L4474 ); 
   and2 U664 ( L3713, L4451, L4476 ); 
   and2 U665 ( L3719, L4451, L4478 ); 
   and2 U666 ( L3725, L4464, L4480 ); 
   and2 U667 ( L3731, L4464, L4482 ); 
   and2 U668 ( L3739, L4464, L4484 ); 
   and2 U669 ( L3745, L4464, L4486 ); 
   and2 U670 ( L3751, L4464, L4488 ); 
   buffer U671 ( L765, L4962 ); 
   buffer U672 ( L765, L5003 ); 
   buffer U673 ( L1007, L5234 ); 
   buffer U674 ( L1007, L5242 ); 
   inv U675 ( L4525, L5250 ); 
   inv U676 ( L579, L5284 ); 
   and2 U677 ( L1488, L2950, L802 ); 
   and2 U678 ( L1482, L2946, L821 ); 
   and2 U679 ( L1477, L2942, L845 ); 
   and2 U680 ( L1471, L2938, L868 ); 
   and2 U681 ( L1464, L2933, L877 ); 
   and2 U682 ( L887, L765, L902 ); 
   or2 U683 ( L777, L907, L908 ); 
   and2 U684 ( L887, L765, L914 ); 
   or2 U685 ( L777, L916, L917 ); 
   and2 U686 ( L887, L765, L953 ); 
   inv U687 ( L1019, L1023 ); 
   and2 U688 ( L1488, L2950, L1035 ); 
   and2 U689 ( L1482, L2946, L1050 ); 
   and2 U690 ( L1477, L2942, L1068 ); 
   and2 U691 ( L1471, L2938, L1086 ); 
   and2 U692 ( L1464, L2933, L1102 ); 
   and2 U693 ( L1019, L1007, L1108 ); 
   or2 U694 ( L1115, L1116, L1117 ); 
   inv U695 ( L5318, L5322 ); 
   and2 U696 ( L1192, L757, L1553 ); 
   and2 U697 ( L1186, L751, L1567 ); 
   and2 U698 ( L2249, L745, L1584 ); 
   and2 U699 ( L2241, L737, L1590 ); 
   and2 U700 ( L1178, L731, L1606 ); 
   and2 U701 ( L2232, L1418, L1624 ); 
   and2 U702 ( L2226, L1412, L1647 ); 
   and2 U703 ( L2220, L1406, L1669 ); 
   and2 U704 ( L2213, L1399, L1677 ); 
   and2 U705 ( L1192, L757, L1802 ); 
   and2 U706 ( L1186, L751, L1816 ); 
   and2 U707 ( L2249, L745, L1834 ); 
   and2 U708 ( L737, L2241, L1841 ); 
   and2 U709 ( L1178, L731, L1866 ); 
   and2 U710 ( L2232, L1418, L1880 ); 
   and2 U711 ( L2226, L1412, L1897 ); 
   and2 U712 ( L2220, L1406, L1914 ); 
   and2 U713 ( L2213, L1399, L1929 ); 
   or2 U714 ( L2045, L2046, L2065 ); 
   or2 U715 ( L2047, L2048, L2069 ); 
   or2 U716 ( L2049, L2050, L2073 ); 
   or2 U717 ( L2051, L2052, L2077 ); 
   or2 U718 ( L2053, L2054, L2081 ); 
   or2 U719 ( L2055, L2056, L2085 ); 
   or2 U720 ( L2057, L2058, L2091 ); 
   or2 U721 ( L2059, L2060, L2099 ); 
   or2 U722 ( L2061, L2062, L2105 ); 
   or2 U723 ( L2063, L2064, L2111 ); 
   or2 U724 ( L2145, L2146, L2163 ); 
   or2 U725 ( L2147, L2148, L2167 ); 
   or2 U726 ( L2149, L2150, L2171 ); 
   or2 U727 ( L2151, L2152, L2175 ); 
   or2 U728 ( L2155, L2156, L2179 ); 
   or2 U729 ( L2157, L2158, L2186 ); 
   or2 U730 ( L2159, L2160, L2192 ); 
   or2 U731 ( L2161, L2162, L2198 ); 
   or2 U732 ( L2297, L2298, L2320 ); 
   or2 U733 ( L2299, L2300, L2323 ); 
   or2 U734 ( L2301, L2302, L2329 ); 
   or2 U735 ( L2303, L2304, L2335 ); 
   and2 U736 ( L4710, L727, L2962 ); 
   and2 U737 ( L4707, L723, L2970 ); 
   and2 U738 ( L4704, L719, L2977 ); 
   and2 U739 ( L4701, L715, L2979 ); 
   and2 U740 ( L4698, L711, L2989 ); 
   and2 U741 ( L4695, L1395, L2998 ); 
   and2 U742 ( L4692, L1391, L3006 ); 
   and2 U743 ( L4689, L1387, L3013 ); 
   and2 U744 ( L4686, L1383, L3015 ); 
   and2 U745 ( L3679, L645, L3183 ); 
   and2 U746 ( L3676, L641, L3192 ); 
   and2 U747 ( L3673, L637, L3200 ); 
   and2 U748 ( L3670, L633, L3207 ); 
   and2 U749 ( L3667, L629, L3209 ); 
   and2 U750 ( L3212, L3170, L3216 ); 
   and2 U751 ( L3170, L3173, L3222 ); 
   inv U752 ( L6690, L6694 ); 
   and2 U753 ( L1535, L2305, L3695 ); 
   or2 U754 ( L3791, L3792, L3816 ); 
   or2 U755 ( L3793, L3794, L3821 ); 
   or2 U756 ( L3795, L3796, L3828 ); 
   or2 U757 ( L3797, L3798, L3833 ); 
   or2 U758 ( L3799, L3800, L3838 ); 
   or2 U759 ( L4125, L4126, L4151 ); 
   or2 U760 ( L4128, L4129, L4154 ); 
   or2 U761 ( L4131, L4132, L4157 ); 
   or2 U762 ( L4134, L4135, L4160 ); 
   or2 U763 ( L4137, L4138, L4163 ); 
   or2 U764 ( L4140, L4141, L4166 ); 
   or2 U765 ( L4143, L4144, L4169 ); 
   or2 U766 ( L4146, L4147, L4172 ); 
   or2 U767 ( L4149, L4150, L4175 ); 
   inv U768 ( L7252, L7256 ); 
   inv U769 ( L7296, L7300 ); 
   or2 U770 ( L4474, L4475, L4490 ); 
   or2 U771 ( L4476, L4477, L4493 ); 
   or2 U772 ( L4478, L4479, L4496 ); 
   or2 U773 ( L4480, L4481, L4499 ); 
   or2 U774 ( L4482, L4483, L4502 ); 
   or2 U775 ( L4484, L4485, L4505 ); 
   or2 U776 ( L4486, L4487, L4508 ); 
   or2 U777 ( L4488, L4489, L4511 ); 
   inv U778 ( L7466, L7470 ); 
   buffer U779 ( L2950, L4884 ); 
   buffer U780 ( L2946, L4892 ); 
   buffer U781 ( L2942, L4900 ); 
   buffer U782 ( L2938, L4908 ); 
   buffer U783 ( L2933, L4924 ); 
   buffer U784 ( L887, L4952 ); 
   nor2 U785 ( L777, L915, L4983 ); 
   buffer U786 ( L887, L4993 ); 
   nor2 U787 ( L1464, L2933, L5011 ); 
   buffer U788 ( L2950, L5194 ); 
   buffer U789 ( L2946, L5202 ); 
   buffer U790 ( L2942, L5210 ); 
   buffer U791 ( L2938, L5218 ); 
   buffer U792 ( L2933, L5226 ); 
   buffer U793 ( L2933, L5247 ); 
   buffer U794 ( L2942, L5255 ); 
   buffer U795 ( L2938, L5258 ); 
   buffer U796 ( L2950, L5263 ); 
   buffer U797 ( L2946, L5266 ); 
   inv U798 ( L5271, L5277 ); 
   inv U799 ( L5274, L5278 ); 
   buffer U800 ( L629, L5281 ); 
   buffer U801 ( L637, L5289 ); 
   buffer U802 ( L633, L5292 ); 
   buffer U803 ( L645, L5297 ); 
   buffer U804 ( L641, L5300 ); 
   inv U805 ( L5305, L5311 ); 
   inv U806 ( L5308, L5312 ); 
   buffer U807 ( L1399, L5315 ); 
   buffer U808 ( L1412, L5323 ); 
   buffer U809 ( L1406, L5326 ); 
   buffer U810 ( L731, L5331 ); 
   buffer U811 ( L1418, L5334 ); 
   buffer U812 ( L745, L5339 ); 
   buffer U813 ( L737, L5342 ); 
   buffer U814 ( L757, L5349 ); 
   buffer U815 ( L751, L5352 ); 
   buffer U816 ( L757, L5396 ); 
   buffer U817 ( L751, L5404 ); 
   buffer U818 ( L745, L5412 ); 
   buffer U819 ( L731, L5420 ); 
   buffer U820 ( L1418, L5428 ); 
   buffer U821 ( L1412, L5436 ); 
   buffer U822 ( L1406, L5444 ); 
   buffer U823 ( L737, L5452 ); 
   buffer U824 ( L1399, L5460 ); 
   nor2 U825 ( L2241, L737, L5465 ); 
   nor2 U826 ( L2213, L1399, L5581 ); 
   buffer U827 ( L757, L5748 ); 
   buffer U828 ( L751, L5756 ); 
   buffer U829 ( L745, L5764 ); 
   buffer U830 ( L737, L5772 ); 
   buffer U831 ( L731, L5780 ); 
   buffer U832 ( L1418, L5788 ); 
   buffer U833 ( L1412, L5796 ); 
   buffer U834 ( L1406, L5804 ); 
   buffer U835 ( L1399, L5812 ); 
   nor2 U836 ( L737, L2241, L5849 ); 
   buffer U837 ( L3682, L5929 ); 
   buffer U838 ( L3682, L6049 ); 
   buffer U839 ( L4710, L6367 ); 
   buffer U840 ( L727, L6370 ); 
   buffer U841 ( L4707, L6375 ); 
   buffer U842 ( L723, L6378 ); 
   buffer U843 ( L4704, L6383 ); 
   buffer U844 ( L719, L6386 ); 
   buffer U845 ( L4698, L6391 ); 
   buffer U846 ( L711, L6394 ); 
   buffer U847 ( L4695, L6399 ); 
   buffer U848 ( L1395, L6402 ); 
   buffer U849 ( L4692, L6407 ); 
   buffer U850 ( L1391, L6410 ); 
   buffer U851 ( L4689, L6415 ); 
   buffer U852 ( L1387, L6418 ); 
   buffer U853 ( L4701, L6423 ); 
   buffer U854 ( L715, L6426 ); 
   buffer U855 ( L4686, L6431 ); 
   buffer U856 ( L1383, L6434 ); 
   buffer U857 ( L3813, L6442 ); 
   buffer U858 ( L3810, L6450 ); 
   buffer U859 ( L3807, L6458 ); 
   buffer U860 ( L3801, L6466 ); 
   buffer U861 ( L3804, L6498 ); 
   buffer U862 ( L3679, L6519 ); 
   buffer U863 ( L645, L6522 ); 
   buffer U864 ( L3676, L6527 ); 
   buffer U865 ( L641, L6530 ); 
   buffer U866 ( L3673, L6535 ); 
   buffer U867 ( L637, L6538 ); 
   buffer U868 ( L3670, L6543 ); 
   buffer U869 ( L633, L6546 ); 
   buffer U870 ( L3667, L6559 ); 
   buffer U871 ( L629, L6562 ); 
   buffer U872 ( L3667, L6687 ); 
   buffer U873 ( L3673, L6695 ); 
   buffer U874 ( L3670, L6698 ); 
   buffer U875 ( L3679, L6703 ); 
   buffer U876 ( L3676, L6706 ); 
   inv U877 ( L6711, L6717 ); 
   inv U878 ( L6714, L6718 ); 
   or2 U879 ( L2153, L2154, L6724 ); 
   or2 U880 ( L2295, L2296, L6768 ); 
   or2 U881 ( L2143, L2144, L7208 ); 
   buffer U882 ( L3801, L7221 ); 
   buffer U883 ( L3807, L7229 ); 
   buffer U884 ( L3804, L7232 ); 
   buffer U885 ( L3813, L7239 ); 
   buffer U886 ( L3810, L7242 ); 
   buffer U887 ( L2305, L7249 ); 
   buffer U888 ( L2312, L7257 ); 
   buffer U889 ( L2308, L7260 ); 
   buffer U890 ( L2316, L7268 ); 
   buffer U891 ( L1383, L7293 ); 
   buffer U892 ( L1391, L7301 ); 
   buffer U893 ( L1387, L7304 ); 
   buffer U894 ( L711, L7309 ); 
   buffer U895 ( L1395, L7312 ); 
   buffer U896 ( L719, L7317 ); 
   buffer U897 ( L715, L7320 ); 
   buffer U898 ( L727, L7327 ); 
   buffer U899 ( L723, L7330 ); 
   buffer U900 ( L2316, L7396 ); 
   buffer U901 ( L2312, L7404 ); 
   buffer U902 ( L2308, L7412 ); 
   buffer U903 ( L3686, L7425 ); 
   buffer U904 ( L4686, L7463 ); 
   buffer U905 ( L4692, L7471 ); 
   buffer U906 ( L4689, L7474 ); 
   buffer U907 ( L4698, L7479 ); 
   buffer U908 ( L4695, L7482 ); 
   buffer U909 ( L4704, L7487 ); 
   buffer U910 ( L4701, L7490 ); 
   buffer U911 ( L4710, L7497 ); 
   buffer U912 ( L4707, L7500 ); 
   or2 U913 ( L4472, L4473, L7507 ); 
   or2 U914 ( L4470, L4471, L7510 ); 
   or2 U915 ( L4122, L4123, L7554 ); 
   nand2 U916 ( L5234, L5237, L1152 ); 
   inv U917 ( L5234, L5238 ); 
   nand2 U918 ( L5242, L5245, L1156 ); 
   inv U919 ( L5242, L5246 ); 
   inv U920 ( L5250, L5254 ); 
   inv U921 ( L5284, L5288 ); 
   or2 U922 ( L3221, L3222, L3223 ); 
   or3 U923 ( L777, L913, L914, L4942 ); 
   inv U924 ( L4962, L4966 ); 
   inv U925 ( L5003, L5007 ); 
   nand2 U926 ( L5274, L5277, L5279 ); 
   nand2 U927 ( L5271, L5278, L5280 ); 
   nand2 U928 ( L5308, L5311, L5313 ); 
   nand2 U929 ( L5305, L5312, L5314 ); 
   nand2 U930 ( L6714, L6717, L6719 ); 
   nand2 U931 ( L6711, L6718, L6720 ); 
   nand2 U932 ( L4884, L4887, L790 ); 
   inv U933 ( L4884, L4888 ); 
   nand2 U934 ( L4892, L4895, L803 ); 
   inv U935 ( L4892, L4896 ); 
   nand2 U936 ( L4900, L4903, L825 ); 
   inv U937 ( L4900, L4904 ); 
   nand2 U938 ( L4908, L4911, L851 ); 
   inv U939 ( L4908, L4912 ); 
   nand2 U940 ( L4924, L4927, L893 ); 
   inv U941 ( L4924, L4928 ); 
   inv U942 ( L902, L906 ); 
   inv U943 ( L908, L912 ); 
   nand2 U944 ( L5194, L5197, L1024 ); 
   inv U945 ( L5194, L5198 ); 
   nand2 U946 ( L5202, L5205, L1036 ); 
   inv U947 ( L5202, L5206 ); 
   nand2 U948 ( L5210, L5213, L1053 ); 
   inv U949 ( L5210, L5214 ); 
   nand2 U950 ( L5218, L5221, L1072 ); 
   inv U951 ( L5218, L5222 ); 
   nand2 U952 ( L5226, L5229, L1091 ); 
   inv U953 ( L5226, L5230 ); 
   inv U954 ( L1108, L1112 ); 
   inv U955 ( L1117, L1121 ); 
   nand2 U956 ( L5231, L5238, L1153 ); 
   nand2 U957 ( L5239, L5246, L1157 ); 
   inv U958 ( L5247, L5253 ); 
   nand2 U959 ( L5247, L5254, L1216 ); 
   inv U960 ( L5255, L5261 ); 
   inv U961 ( L5258, L5262 ); 
   inv U962 ( L5263, L5269 ); 
   inv U963 ( L5266, L5270 ); 
   inv U964 ( L5281, L5287 ); 
   nand2 U965 ( L5281, L5288, L1239 ); 
   inv U966 ( L5289, L5295 ); 
   inv U967 ( L5292, L5296 ); 
   inv U968 ( L5297, L5303 ); 
   inv U969 ( L5300, L5304 ); 
   inv U970 ( L5315, L5321 ); 
   nand2 U971 ( L5315, L5322, L1262 ); 
   inv U972 ( L5323, L5329 ); 
   inv U973 ( L5326, L5330 ); 
   inv U974 ( L5331, L5337 ); 
   inv U975 ( L5334, L5338 ); 
   nand2 U976 ( L5396, L5399, L1544 ); 
   inv U977 ( L5396, L5400 ); 
   nand2 U978 ( L5404, L5407, L1554 ); 
   inv U979 ( L5404, L5408 ); 
   nand2 U980 ( L5412, L5415, L1571 ); 
   inv U981 ( L5412, L5416 ); 
   nand2 U982 ( L5420, L5423, L1596 ); 
   inv U983 ( L5420, L5424 ); 
   nand2 U984 ( L5428, L5431, L1607 ); 
   inv U985 ( L5428, L5432 ); 
   nand2 U986 ( L5436, L5439, L1628 ); 
   inv U987 ( L5436, L5440 ); 
   nand2 U988 ( L5444, L5447, L1653 ); 
   inv U989 ( L5444, L5448 ); 
   nand2 U990 ( L5452, L5455, L1685 ); 
   inv U991 ( L5452, L5456 ); 
   nand2 U992 ( L5460, L5463, L1693 ); 
   inv U993 ( L5460, L5464 ); 
   nand2 U994 ( L5748, L5751, L1793 ); 
   inv U995 ( L5748, L5752 ); 
   nand2 U996 ( L5756, L5759, L1803 ); 
   inv U997 ( L5756, L5760 ); 
   nand2 U998 ( L5764, L5767, L1820 ); 
   inv U999 ( L5764, L5768 ); 
   nand2 U1000 ( L5772, L5775, L1848 ); 
   inv U1001 ( L5772, L5776 ); 
   nand2 U1002 ( L5780, L5783, L1857 ); 
   inv U1003 ( L5780, L5784 ); 
   nand2 U1004 ( L5788, L5791, L1867 ); 
   inv U1005 ( L5788, L5792 ); 
   nand2 U1006 ( L5796, L5799, L1883 ); 
   inv U1007 ( L5796, L5800 ); 
   nand2 U1008 ( L5804, L5807, L1901 ); 
   inv U1009 ( L5804, L5808 ); 
   nand2 U1010 ( L5812, L5815, L1919 ); 
   inv U1011 ( L5812, L5816 ); 
   inv U1012 ( L5849, L5855 ); 
   and2 U1013 ( L3751, L2111, L2351 ); 
   and2 U1014 ( L3745, L2105, L2366 ); 
   and2 U1015 ( L3739, L2099, L2384 ); 
   and2 U1016 ( L2091, L3731, L2391 ); 
   and2 U1017 ( L3725, L2085, L2417 ); 
   and2 U1018 ( L3719, L2335, L2431 ); 
   and2 U1019 ( L3713, L2329, L2448 ); 
   and2 U1020 ( L3707, L2323, L2465 ); 
   inv U1021 ( L5929, L5935 ); 
   and2 U1022 ( L3751, L2111, L2597 ); 
   and2 U1023 ( L3745, L2105, L2612 ); 
   and2 U1024 ( L3739, L2099, L2629 ); 
   and2 U1025 ( L3731, L2091, L2635 ); 
   and2 U1026 ( L3725, L2085, L2652 ); 
   and2 U1027 ( L3719, L2335, L2670 ); 
   and2 U1028 ( L3713, L2329, L2693 ); 
   and2 U1029 ( L3707, L2323, L2715 ); 
   inv U1030 ( L6049, L6055 ); 
   inv U1031 ( L6367, L6373 ); 
   inv U1032 ( L6370, L6374 ); 
   inv U1033 ( L6375, L6381 ); 
   inv U1034 ( L6378, L6382 ); 
   inv U1035 ( L6383, L6389 ); 
   inv U1036 ( L6386, L6390 ); 
   inv U1037 ( L6391, L6397 ); 
   inv U1038 ( L6394, L6398 ); 
   inv U1039 ( L6399, L6405 ); 
   inv U1040 ( L6402, L6406 ); 
   inv U1041 ( L6407, L6413 ); 
   inv U1042 ( L6410, L6414 ); 
   inv U1043 ( L6415, L6421 ); 
   inv U1044 ( L6418, L6422 ); 
   inv U1045 ( L6423, L6429 ); 
   inv U1046 ( L6426, L6430 ); 
   inv U1047 ( L6431, L6437 ); 
   inv U1048 ( L6434, L6438 ); 
   inv U1049 ( L6442, L6446 ); 
   and2 U1050 ( L4175, L3813, L3059 ); 
   inv U1051 ( L6450, L6454 ); 
   and2 U1052 ( L4172, L3810, L3068 ); 
   inv U1053 ( L6458, L6462 ); 
   and2 U1054 ( L4169, L3807, L3076 ); 
   and2 U1055 ( L4166, L3804, L3079 ); 
   inv U1056 ( L6466, L6470 ); 
   and2 U1057 ( L4163, L3801, L3090 ); 
   and2 U1058 ( L4160, L2175, L3099 ); 
   and2 U1059 ( L4157, L2171, L3107 ); 
   and2 U1060 ( L4154, L2167, L3114 ); 
   and2 U1061 ( L4151, L2163, L3116 ); 
   inv U1062 ( L6498, L6502 ); 
   inv U1063 ( L6519, L6525 ); 
   inv U1064 ( L6522, L6526 ); 
   inv U1065 ( L6527, L6533 ); 
   inv U1066 ( L6530, L6534 ); 
   inv U1067 ( L6535, L6541 ); 
   inv U1068 ( L6538, L6542 ); 
   inv U1069 ( L6543, L6549 ); 
   inv U1070 ( L6546, L6550 ); 
   inv U1071 ( L6559, L6565 ); 
   inv U1072 ( L6562, L6566 ); 
   inv U1073 ( L3216, L3220 ); 
   and2 U1074 ( L4439, L3838, L3292 ); 
   and2 U1075 ( L4434, L3833, L3308 ); 
   and2 U1076 ( L4429, L3828, L3327 ); 
   and2 U1077 ( L3821, L4422, L3335 ); 
   and2 U1078 ( L4417, L3816, L3362 ); 
   and2 U1079 ( L4412, L2198, L3376 ); 
   and2 U1080 ( L4407, L2192, L3393 ); 
   and2 U1081 ( L4402, L2186, L3410 ); 
   and2 U1082 ( L4396, L2179, L3425 ); 
   inv U1083 ( L6687, L6693 ); 
   nand2 U1084 ( L6687, L6694, L3503 ); 
   inv U1085 ( L6695, L6701 ); 
   inv U1086 ( L6698, L6702 ); 
   inv U1087 ( L6703, L6709 ); 
   inv U1088 ( L6706, L6710 ); 
   inv U1089 ( L6724, L6728 ); 
   inv U1090 ( L6768, L6772 ); 
   and2 U1091 ( L4439, L3838, L3853 ); 
   and2 U1092 ( L4434, L3833, L3868 ); 
   and2 U1093 ( L4429, L3828, L3885 ); 
   and2 U1094 ( L4422, L3821, L3891 ); 
   and2 U1095 ( L4417, L3816, L3908 ); 
   and2 U1096 ( L4412, L2198, L3926 ); 
   and2 U1097 ( L4407, L2192, L3949 ); 
   and2 U1098 ( L4402, L2186, L3971 ); 
   and2 U1099 ( L4396, L2179, L3979 ); 
   inv U1100 ( L7208, L7212 ); 
   inv U1101 ( L7221, L7227 ); 
   inv U1102 ( L7249, L7255 ); 
   nand2 U1103 ( L7249, L7256, L4202 ); 
   inv U1104 ( L7257, L7263 ); 
   inv U1105 ( L7260, L7264 ); 
   inv U1106 ( L7268, L7272 ); 
   inv U1107 ( L7293, L7299 ); 
   nand2 U1108 ( L7293, L7300, L4225 ); 
   inv U1109 ( L7301, L7307 ); 
   inv U1110 ( L7304, L7308 ); 
   inv U1111 ( L7309, L7315 ); 
   inv U1112 ( L7312, L7316 ); 
   and2 U1113 ( L4511, L2081, L4297 ); 
   and2 U1114 ( L4508, L2077, L4305 ); 
   and2 U1115 ( L4505, L2073, L4312 ); 
   and2 U1116 ( L4502, L2069, L4314 ); 
   and2 U1117 ( L4499, L2065, L4324 ); 
   inv U1118 ( L7396, L7400 ); 
   and2 U1119 ( L4496, L2316, L4333 ); 
   inv U1120 ( L7404, L7408 ); 
   and2 U1121 ( L4493, L2312, L4341 ); 
   inv U1122 ( L7412, L7416 ); 
   and2 U1123 ( L4490, L2308, L4348 ); 
   and2 U1124 ( L3686, L3695, L4349 ); 
   inv U1125 ( L7425, L7431 ); 
   and2 U1126 ( L2320, L1535, L4389 ); 
   inv U1127 ( L7463, L7469 ); 
   nand2 U1128 ( L7463, L7470, L4530 ); 
   inv U1129 ( L7471, L7477 ); 
   inv U1130 ( L7474, L7478 ); 
   inv U1131 ( L7479, L7485 ); 
   inv U1132 ( L7482, L7486 ); 
   inv U1133 ( L7507, L7513 ); 
   inv U1134 ( L7510, L7514 ); 
   inv U1135 ( L7554, L7558 ); 
   or2 U1136 ( L917, L953, L4932 ); 
   inv U1137 ( L4952, L4956 ); 
   inv U1138 ( L917, L4973 ); 
   inv U1139 ( L4983, L4987 ); 
   inv U1140 ( L4993, L4997 ); 
   inv U1141 ( L5011, L5017 ); 
   buffer U1142 ( L877, L5099 ); 
   inv U1143 ( L5339, L5345 ); 
   inv U1144 ( L5342, L5346 ); 
   inv U1145 ( L5349, L5355 ); 
   inv U1146 ( L5352, L5356 ); 
   nand2 U1147 ( L5279, L5280, L5372 ); 
   nand2 U1148 ( L5313, L5314, L5380 ); 
   inv U1149 ( L5465, L5471 ); 
   buffer U1150 ( L1590, L5523 ); 
   inv U1151 ( L5581, L5587 ); 
   buffer U1152 ( L1677, L5669 ); 
   buffer U1153 ( L1841, L5857 ); 
   buffer U1154 ( L2111, L5868 ); 
   buffer U1155 ( L2105, L5876 ); 
   buffer U1156 ( L2099, L5884 ); 
   buffer U1157 ( L2091, L5892 ); 
   buffer U1158 ( L2085, L5900 ); 
   buffer U1159 ( L2335, L5908 ); 
   buffer U1160 ( L2329, L5916 ); 
   buffer U1161 ( L2323, L5924 ); 
   nor2 U1162 ( L2091, L3731, L5969 ); 
   buffer U1163 ( L2111, L5988 ); 
   buffer U1164 ( L2105, L5996 ); 
   buffer U1165 ( L2099, L6004 ); 
   buffer U1166 ( L2085, L6012 ); 
   buffer U1167 ( L2335, L6020 ); 
   buffer U1168 ( L2329, L6028 ); 
   buffer U1169 ( L2323, L6036 ); 
   buffer U1170 ( L2091, L6044 ); 
   nor2 U1171 ( L3731, L2091, L6057 ); 
   buffer U1172 ( L4175, L6439 ); 
   buffer U1173 ( L4172, L6447 ); 
   buffer U1174 ( L4169, L6455 ); 
   buffer U1175 ( L4163, L6463 ); 
   buffer U1176 ( L4160, L6471 ); 
   buffer U1177 ( L2175, L6474 ); 
   buffer U1178 ( L4157, L6479 ); 
   buffer U1179 ( L2171, L6482 ); 
   buffer U1180 ( L4154, L6487 ); 
   buffer U1181 ( L2167, L6490 ); 
   buffer U1182 ( L4166, L6495 ); 
   buffer U1183 ( L4151, L6503 ); 
   buffer U1184 ( L2163, L6506 ); 
   buffer U1185 ( L3838, L6570 ); 
   buffer U1186 ( L3833, L6578 ); 
   buffer U1187 ( L3828, L6586 ); 
   buffer U1188 ( L3821, L6594 ); 
   buffer U1189 ( L3816, L6602 ); 
   buffer U1190 ( L2198, L6610 ); 
   buffer U1191 ( L2192, L6618 ); 
   buffer U1192 ( L2186, L6626 ); 
   buffer U1193 ( L2179, L6634 ); 
   nor2 U1194 ( L3821, L4422, L6671 ); 
   buffer U1195 ( L2179, L6721 ); 
   buffer U1196 ( L2192, L6729 ); 
   buffer U1197 ( L2186, L6732 ); 
   buffer U1198 ( L3816, L6737 ); 
   buffer U1199 ( L2198, L6740 ); 
   buffer U1200 ( L3828, L6745 ); 
   buffer U1201 ( L3821, L6748 ); 
   buffer U1202 ( L3838, L6755 ); 
   buffer U1203 ( L3833, L6758 ); 
   buffer U1204 ( L2320, L6765 ); 
   buffer U1205 ( L2329, L6773 ); 
   buffer U1206 ( L2323, L6776 ); 
   buffer U1207 ( L2085, L6781 ); 
   buffer U1208 ( L2335, L6784 ); 
   buffer U1209 ( L2099, L6789 ); 
   buffer U1210 ( L2091, L6792 ); 
   buffer U1211 ( L2111, L6799 ); 
   buffer U1212 ( L2105, L6802 ); 
   nand2 U1213 ( L6719, L6720, L6832 ); 
   buffer U1214 ( L3838, L6856 ); 
   buffer U1215 ( L3833, L6864 ); 
   buffer U1216 ( L3828, L6872 ); 
   buffer U1217 ( L3816, L6880 ); 
   buffer U1218 ( L2198, L6888 ); 
   buffer U1219 ( L2192, L6896 ); 
   buffer U1220 ( L2186, L6904 ); 
   buffer U1221 ( L3821, L6912 ); 
   buffer U1222 ( L2179, L6920 ); 
   nor2 U1223 ( L4422, L3821, L6925 ); 
   nor2 U1224 ( L4396, L2179, L7041 ); 
   buffer U1225 ( L2163, L7205 ); 
   buffer U1226 ( L2171, L7213 ); 
   buffer U1227 ( L2167, L7216 ); 
   buffer U1228 ( L2175, L7224 ); 
   inv U1229 ( L7229, L7235 ); 
   inv U1230 ( L7232, L7236 ); 
   inv U1231 ( L7239, L7245 ); 
   inv U1232 ( L7242, L7246 ); 
   buffer U1233 ( L2065, L7265 ); 
   buffer U1234 ( L2073, L7273 ); 
   buffer U1235 ( L2069, L7276 ); 
   buffer U1236 ( L2081, L7283 ); 
   buffer U1237 ( L2077, L7286 ); 
   inv U1238 ( L7317, L7323 ); 
   inv U1239 ( L7320, L7324 ); 
   inv U1240 ( L7327, L7333 ); 
   inv U1241 ( L7330, L7334 ); 
   buffer U1242 ( L4511, L7361 ); 
   buffer U1243 ( L2081, L7364 ); 
   buffer U1244 ( L4508, L7369 ); 
   buffer U1245 ( L2077, L7372 ); 
   buffer U1246 ( L4505, L7377 ); 
   buffer U1247 ( L2073, L7380 ); 
   buffer U1248 ( L4499, L7385 ); 
   buffer U1249 ( L2065, L7388 ); 
   buffer U1250 ( L4496, L7393 ); 
   buffer U1251 ( L4493, L7401 ); 
   buffer U1252 ( L4490, L7409 ); 
   buffer U1253 ( L4502, L7417 ); 
   buffer U1254 ( L2069, L7420 ); 
   buffer U1255 ( L3695, L7428 ); 
   inv U1256 ( L7487, L7493 ); 
   inv U1257 ( L7490, L7494 ); 
   inv U1258 ( L7497, L7503 ); 
   inv U1259 ( L7500, L7504 ); 
   buffer U1260 ( L4493, L7515 ); 
   buffer U1261 ( L4490, L7518 ); 
   buffer U1262 ( L4499, L7523 ); 
   buffer U1263 ( L4496, L7526 ); 
   buffer U1264 ( L4505, L7531 ); 
   buffer U1265 ( L4502, L7534 ); 
   buffer U1266 ( L4511, L7541 ); 
   buffer U1267 ( L4508, L7544 ); 
   buffer U1268 ( L4151, L7551 ); 
   buffer U1269 ( L4157, L7559 ); 
   buffer U1270 ( L4154, L7562 ); 
   buffer U1271 ( L4163, L7567 ); 
   buffer U1272 ( L4160, L7570 ); 
   buffer U1273 ( L4169, L7575 ); 
   buffer U1274 ( L4166, L7578 ); 
   buffer U1275 ( L4175, L7585 ); 
   buffer U1276 ( L4172, L7588 ); 
   nand2 U1277 ( L1121, L1112, L1176 ); 
   nand2 U1278 ( L912, L906, L957 ); 
   nand2 U1279 ( L4881, L4888, L791 ); 
   nand2 U1280 ( L4889, L4896, L804 ); 
   nand2 U1281 ( L4897, L4904, L826 ); 
   nand2 U1282 ( L4905, L4912, L852 ); 
   nand2 U1283 ( L4921, L4928, L894 ); 
   nand2 U1284 ( L5191, L5198, L1025 ); 
   nand2 U1285 ( L5199, L5206, L1037 ); 
   nand2 U1286 ( L5207, L5214, L1054 ); 
   nand2 U1287 ( L5215, L5222, L1073 ); 
   nand2 U1288 ( L5223, L5230, L1092 ); 
   nand2 U1289 ( L1152, L1153, L1154 ); 
   nand2 U1290 ( L1156, L1157, L1158 ); 
   nand2 U1291 ( L5250, L5253, L1215 ); 
   nand2 U1292 ( L5258, L5261, L1224 ); 
   nand2 U1293 ( L5255, L5262, L1225 ); 
   nand2 U1294 ( L5266, L5269, L1233 ); 
   nand2 U1295 ( L5263, L5270, L1234 ); 
   nand2 U1296 ( L5284, L5287, L1238 ); 
   nand2 U1297 ( L5292, L5295, L1247 ); 
   nand2 U1298 ( L5289, L5296, L1248 ); 
   nand2 U1299 ( L5300, L5303, L1256 ); 
   nand2 U1300 ( L5297, L5304, L1257 ); 
   nand2 U1301 ( L5318, L5321, L1261 ); 
   nand2 U1302 ( L5326, L5329, L1270 ); 
   nand2 U1303 ( L5323, L5330, L1271 ); 
   nand2 U1304 ( L5334, L5337, L1279 ); 
   nand2 U1305 ( L5331, L5338, L1280 ); 
   nand2 U1306 ( L5393, L5400, L1545 ); 
   nand2 U1307 ( L5401, L5408, L1555 ); 
   nand2 U1308 ( L5409, L5416, L1572 ); 
   nand2 U1309 ( L5417, L5424, L1597 ); 
   nand2 U1310 ( L5425, L5432, L1608 ); 
   nand2 U1311 ( L5433, L5440, L1629 ); 
   nand2 U1312 ( L5441, L5448, L1654 ); 
   nand2 U1313 ( L5449, L5456, L1686 ); 
   nand2 U1314 ( L5457, L5464, L1694 ); 
   nand2 U1315 ( L5745, L5752, L1794 ); 
   nand2 U1316 ( L5753, L5760, L1804 ); 
   nand2 U1317 ( L5761, L5768, L1821 ); 
   nand2 U1318 ( L5769, L5776, L1849 ); 
   nand2 U1319 ( L5777, L5784, L1858 ); 
   nand2 U1320 ( L5785, L5792, L1868 ); 
   nand2 U1321 ( L5793, L5800, L1884 ); 
   nand2 U1322 ( L5801, L5808, L1902 ); 
   nand2 U1323 ( L5809, L5816, L1920 ); 
   nand2 U1324 ( L6370, L6373, L2954 ); 
   nand2 U1325 ( L6367, L6374, L2955 ); 
   nand2 U1326 ( L6378, L6381, L2963 ); 
   nand2 U1327 ( L6375, L6382, L2964 ); 
   nand2 U1328 ( L6386, L6389, L2971 ); 
   nand2 U1329 ( L6383, L6390, L2972 ); 
   nand2 U1330 ( L6394, L6397, L2980 ); 
   nand2 U1331 ( L6391, L6398, L2981 ); 
   nand2 U1332 ( L6402, L6405, L2990 ); 
   nand2 U1333 ( L6399, L6406, L2991 ); 
   nand2 U1334 ( L6410, L6413, L2999 ); 
   nand2 U1335 ( L6407, L6414, L3000 ); 
   nand2 U1336 ( L6418, L6421, L3007 ); 
   nand2 U1337 ( L6415, L6422, L3008 ); 
   nand2 U1338 ( L6426, L6429, L3016 ); 
   nand2 U1339 ( L6423, L6430, L3017 ); 
   nand2 U1340 ( L6434, L6437, L3019 ); 
   nand2 U1341 ( L6431, L6438, L3020 ); 
   nand2 U1342 ( L6522, L6525, L3174 ); 
   nand2 U1343 ( L6519, L6526, L3175 ); 
   nand2 U1344 ( L6530, L6533, L3184 ); 
   nand2 U1345 ( L6527, L6534, L3185 ); 
   nand2 U1346 ( L6538, L6541, L3193 ); 
   nand2 U1347 ( L6535, L6542, L3194 ); 
   nand2 U1348 ( L6546, L6549, L3201 ); 
   nand2 U1349 ( L6543, L6550, L3202 ); 
   nand2 U1350 ( L6562, L6565, L3213 ); 
   nand2 U1351 ( L6559, L6566, L3214 ); 
   inv U1352 ( L3223, L3227 ); 
   nand2 U1353 ( L6690, L6693, L3502 ); 
   nand2 U1354 ( L6698, L6701, L3511 ); 
   nand2 U1355 ( L6695, L6702, L3512 ); 
   nand2 U1356 ( L6706, L6709, L3520 ); 
   nand2 U1357 ( L6703, L6710, L3521 ); 
   nand2 U1358 ( L7252, L7255, L4201 ); 
   nand2 U1359 ( L7260, L7263, L4210 ); 
   nand2 U1360 ( L7257, L7264, L4211 ); 
   nand2 U1361 ( L7296, L7299, L4224 ); 
   nand2 U1362 ( L7304, L7307, L4233 ); 
   nand2 U1363 ( L7301, L7308, L4234 ); 
   nand2 U1364 ( L7312, L7315, L4242 ); 
   nand2 U1365 ( L7309, L7316, L4243 ); 
   nand2 U1366 ( L7466, L7469, L4529 ); 
   nand2 U1367 ( L7474, L7477, L4538 ); 
   nand2 U1368 ( L7471, L7478, L4539 ); 
   nand2 U1369 ( L7482, L7485, L4547 ); 
   nand2 U1370 ( L7479, L7486, L4548 ); 
   nand2 U1371 ( L7510, L7513, L4552 ); 
   nand2 U1372 ( L7507, L7514, L4553 ); 
   inv U1373 ( L4942, L4946 ); 
   nand2 U1374 ( L5342, L5345, L5347 ); 
   nand2 U1375 ( L5339, L5346, L5348 ); 
   nand2 U1376 ( L5352, L5355, L5357 ); 
   nand2 U1377 ( L5349, L5356, L5358 ); 
   nand2 U1378 ( L7232, L7235, L7237 ); 
   nand2 U1379 ( L7229, L7236, L7238 ); 
   nand2 U1380 ( L7242, L7245, L7247 ); 
   nand2 U1381 ( L7239, L7246, L7248 ); 
   nand2 U1382 ( L7320, L7323, L7325 ); 
   nand2 U1383 ( L7317, L7324, L7326 ); 
   nand2 U1384 ( L7330, L7333, L7335 ); 
   nand2 U1385 ( L7327, L7334, L7336 ); 
   nand2 U1386 ( L7490, L7493, L7495 ); 
   nand2 U1387 ( L7487, L7494, L7496 ); 
   nand2 U1388 ( L7500, L7503, L7505 ); 
   nand2 U1389 ( L7497, L7504, L7506 ); 
   nand2 U1390 ( L3227, L3220, L3244 ); 
   nand2 U1391 ( L790, L791, L792 ); 
   nand2 U1392 ( L803, L804, L805 ); 
   nand2 U1393 ( L825, L826, L827 ); 
   nand2 U1394 ( L851, L852, L853 ); 
   nand2 U1395 ( L893, L894, L895 ); 
   nand2 U1396 ( L1024, L1025, L1026 ); 
   nand2 U1397 ( L1036, L1037, L1038 ); 
   nand2 U1398 ( L1053, L1054, L1055 ); 
   nand2 U1399 ( L1072, L1073, L1074 ); 
   nand2 U1400 ( L1091, L1092, L1093 ); 
   inv U1401 ( L1154, L1155 ); 
   nand2 U1402 ( L1215, L1216, L1217 ); 
   nand2 U1403 ( L1224, L1225, L1226 ); 
   nand2 U1404 ( L1233, L1234, L1235 ); 
   nand2 U1405 ( L1238, L1239, L1240 ); 
   nand2 U1406 ( L1247, L1248, L1249 ); 
   nand2 U1407 ( L1256, L1257, L1258 ); 
   nand2 U1408 ( L1261, L1262, L1263 ); 
   nand2 U1409 ( L1270, L1271, L1272 ); 
   nand2 U1410 ( L1279, L1280, L1281 ); 
   inv U1411 ( L5372, L5376 ); 
   inv U1412 ( L5380, L5384 ); 
   nand2 U1413 ( L1544, L1545, L1546 ); 
   nand2 U1414 ( L1554, L1555, L1556 ); 
   nand2 U1415 ( L1571, L1572, L1573 ); 
   nand2 U1416 ( L1596, L1597, L1598 ); 
   nand2 U1417 ( L1607, L1608, L1609 ); 
   nand2 U1418 ( L1628, L1629, L1630 ); 
   nand2 U1419 ( L1653, L1654, L1655 ); 
   nand2 U1420 ( L1685, L1686, L1687 ); 
   nand2 U1421 ( L1693, L1694, L1695 ); 
   nand2 U1422 ( L1793, L1794, L1795 ); 
   nand2 U1423 ( L1803, L1804, L1805 ); 
   nand2 U1424 ( L1820, L1821, L1822 ); 
   nand2 U1425 ( L1848, L1849, L1850 ); 
   nand2 U1426 ( L1857, L1858, L1859 ); 
   nand2 U1427 ( L1867, L1868, L1869 ); 
   nand2 U1428 ( L1883, L1884, L1885 ); 
   nand2 U1429 ( L1901, L1902, L1903 ); 
   nand2 U1430 ( L1919, L1920, L1921 ); 
   inv U1431 ( L5857, L5863 ); 
   nand2 U1432 ( L5868, L5871, L2341 ); 
   inv U1433 ( L5868, L5872 ); 
   nand2 U1434 ( L5876, L5879, L2352 ); 
   inv U1435 ( L5876, L5880 ); 
   nand2 U1436 ( L5884, L5887, L2370 ); 
   inv U1437 ( L5884, L5888 ); 
   nand2 U1438 ( L5892, L5895, L2398 ); 
   inv U1439 ( L5892, L5896 ); 
   nand2 U1440 ( L5900, L5903, L2407 ); 
   inv U1441 ( L5900, L5904 ); 
   nand2 U1442 ( L5908, L5911, L2418 ); 
   inv U1443 ( L5908, L5912 ); 
   nand2 U1444 ( L5916, L5919, L2434 ); 
   inv U1445 ( L5916, L5920 ); 
   nand2 U1446 ( L5924, L5927, L2452 ); 
   inv U1447 ( L5924, L5928 ); 
   and2 U1448 ( L3682, L4389, L2481 ); 
   inv U1449 ( L5969, L5975 ); 
   nand2 U1450 ( L5988, L5991, L2587 ); 
   inv U1451 ( L5988, L5992 ); 
   nand2 U1452 ( L5996, L5999, L2598 ); 
   inv U1453 ( L5996, L6000 ); 
   nand2 U1454 ( L6004, L6007, L2616 ); 
   inv U1455 ( L6004, L6008 ); 
   nand2 U1456 ( L6012, L6015, L2641 ); 
   inv U1457 ( L6012, L6016 ); 
   nand2 U1458 ( L6020, L6023, L2653 ); 
   inv U1459 ( L6020, L6024 ); 
   nand2 U1460 ( L6028, L6031, L2674 ); 
   inv U1461 ( L6028, L6032 ); 
   nand2 U1462 ( L6036, L6039, L2699 ); 
   inv U1463 ( L6036, L6040 ); 
   and2 U1464 ( L3682, L4389, L2724 ); 
   nand2 U1465 ( L6044, L6047, L2732 ); 
   inv U1466 ( L6044, L6048 ); 
   nand2 U1467 ( L2954, L2955, L2956 ); 
   nand2 U1468 ( L2963, L2964, L2965 ); 
   nand2 U1469 ( L2971, L2972, L2973 ); 
   nand2 U1470 ( L2980, L2981, L2982 ); 
   nand2 U1471 ( L2990, L2991, L2992 ); 
   nand2 U1472 ( L2999, L3000, L3001 ); 
   nand2 U1473 ( L3007, L3008, L3009 ); 
   nand2 U1474 ( L3016, L3017, L3018 ); 
   nand2 U1475 ( L3019, L3020, L3021 ); 
   inv U1476 ( L6439, L6445 ); 
   nand2 U1477 ( L6439, L6446, L3051 ); 
   inv U1478 ( L6447, L6453 ); 
   nand2 U1479 ( L6447, L6454, L3061 ); 
   inv U1480 ( L6455, L6461 ); 
   nand2 U1481 ( L6455, L6462, L3070 ); 
   inv U1482 ( L6463, L6469 ); 
   nand2 U1483 ( L6463, L6470, L3081 ); 
   inv U1484 ( L6471, L6477 ); 
   inv U1485 ( L6474, L6478 ); 
   inv U1486 ( L6479, L6485 ); 
   inv U1487 ( L6482, L6486 ); 
   inv U1488 ( L6487, L6493 ); 
   inv U1489 ( L6490, L6494 ); 
   inv U1490 ( L6495, L6501 ); 
   nand2 U1491 ( L6495, L6502, L3118 ); 
   inv U1492 ( L6503, L6509 ); 
   inv U1493 ( L6506, L6510 ); 
   nand2 U1494 ( L3174, L3175, L3176 ); 
   nand2 U1495 ( L3184, L3185, L3186 ); 
   nand2 U1496 ( L3193, L3194, L3195 ); 
   nand2 U1497 ( L3201, L3202, L3203 ); 
   nand2 U1498 ( L3213, L3214, L3215 ); 
   nand2 U1499 ( L6570, L6573, L3281 ); 
   inv U1500 ( L6570, L6574 ); 
   nand2 U1501 ( L6578, L6581, L3293 ); 
   inv U1502 ( L6578, L6582 ); 
   nand2 U1503 ( L6586, L6589, L3312 ); 
   inv U1504 ( L6586, L6590 ); 
   nand2 U1505 ( L6594, L6597, L3342 ); 
   inv U1506 ( L6594, L6598 ); 
   nand2 U1507 ( L6602, L6605, L3351 ); 
   inv U1508 ( L6602, L6606 ); 
   nand2 U1509 ( L6610, L6613, L3363 ); 
   inv U1510 ( L6610, L6614 ); 
   nand2 U1511 ( L6618, L6621, L3379 ); 
   inv U1512 ( L6618, L6622 ); 
   nand2 U1513 ( L6626, L6629, L3397 ); 
   inv U1514 ( L6626, L6630 ); 
   nand2 U1515 ( L6634, L6637, L3415 ); 
   inv U1516 ( L6634, L6638 ); 
   inv U1517 ( L6671, L6677 ); 
   nand2 U1518 ( L3502, L3503, L3504 ); 
   nand2 U1519 ( L3511, L3512, L3513 ); 
   nand2 U1520 ( L3520, L3521, L3522 ); 
   inv U1521 ( L6721, L6727 ); 
   nand2 U1522 ( L6721, L6728, L3526 ); 
   inv U1523 ( L6729, L6735 ); 
   inv U1524 ( L6732, L6736 ); 
   inv U1525 ( L6737, L6743 ); 
   inv U1526 ( L6740, L6744 ); 
   inv U1527 ( L6765, L6771 ); 
   nand2 U1528 ( L6765, L6772, L3549 ); 
   inv U1529 ( L6773, L6779 ); 
   inv U1530 ( L6776, L6780 ); 
   inv U1531 ( L6781, L6787 ); 
   inv U1532 ( L6784, L6788 ); 
   inv U1533 ( L6832, L6836 ); 
   nand2 U1534 ( L6856, L6859, L3843 ); 
   inv U1535 ( L6856, L6860 ); 
   nand2 U1536 ( L6864, L6867, L3854 ); 
   inv U1537 ( L6864, L6868 ); 
   nand2 U1538 ( L6872, L6875, L3872 ); 
   inv U1539 ( L6872, L6876 ); 
   nand2 U1540 ( L6880, L6883, L3897 ); 
   inv U1541 ( L6880, L6884 ); 
   nand2 U1542 ( L6888, L6891, L3909 ); 
   inv U1543 ( L6888, L6892 ); 
   nand2 U1544 ( L6896, L6899, L3930 ); 
   inv U1545 ( L6896, L6900 ); 
   nand2 U1546 ( L6904, L6907, L3955 ); 
   inv U1547 ( L6904, L6908 ); 
   nand2 U1548 ( L6912, L6915, L3987 ); 
   inv U1549 ( L6912, L6916 ); 
   nand2 U1550 ( L6920, L6923, L3995 ); 
   inv U1551 ( L6920, L6924 ); 
   inv U1552 ( L7205, L7211 ); 
   nand2 U1553 ( L7205, L7212, L4179 ); 
   inv U1554 ( L7213, L7219 ); 
   inv U1555 ( L7216, L7220 ); 
   nand2 U1556 ( L7224, L7227, L4196 ); 
   inv U1557 ( L7224, L7228 ); 
   nand2 U1558 ( L4201, L4202, L4203 ); 
   nand2 U1559 ( L4210, L4211, L4212 ); 
   inv U1560 ( L7265, L7271 ); 
   nand2 U1561 ( L7265, L7272, L4220 ); 
   nand2 U1562 ( L4224, L4225, L4226 ); 
   nand2 U1563 ( L4233, L4234, L4235 ); 
   nand2 U1564 ( L4242, L4243, L4244 ); 
   inv U1565 ( L7361, L7367 ); 
   inv U1566 ( L7364, L7368 ); 
   inv U1567 ( L7369, L7375 ); 
   inv U1568 ( L7372, L7376 ); 
   inv U1569 ( L7377, L7383 ); 
   inv U1570 ( L7380, L7384 ); 
   inv U1571 ( L7385, L7391 ); 
   inv U1572 ( L7388, L7392 ); 
   inv U1573 ( L7393, L7399 ); 
   nand2 U1574 ( L7393, L7400, L4326 ); 
   inv U1575 ( L7401, L7407 ); 
   nand2 U1576 ( L7401, L7408, L4335 ); 
   inv U1577 ( L7409, L7415 ); 
   nand2 U1578 ( L7409, L7416, L4343 ); 
   inv U1579 ( L7417, L7423 ); 
   inv U1580 ( L7420, L7424 ); 
   nand2 U1581 ( L7428, L7431, L4353 ); 
   inv U1582 ( L7428, L7432 ); 
   nand2 U1583 ( L4529, L4530, L4531 ); 
   nand2 U1584 ( L4538, L4539, L4540 ); 
   nand2 U1585 ( L4547, L4548, L4549 ); 
   nand2 U1586 ( L4552, L4553, L4554 ); 
   inv U1587 ( L7515, L7521 ); 
   inv U1588 ( L7518, L7522 ); 
   inv U1589 ( L7523, L7529 ); 
   inv U1590 ( L7526, L7530 ); 
   inv U1591 ( L7551, L7557 ); 
   nand2 U1592 ( L7551, L7558, L4576 ); 
   inv U1593 ( L7559, L7565 ); 
   inv U1594 ( L7562, L7566 ); 
   inv U1595 ( L7567, L7573 ); 
   inv U1596 ( L7570, L7574 ); 
   inv U1597 ( L4932, L4936 ); 
   nand2 U1598 ( L4932, L4935, L4937 ); 
   inv U1599 ( L4973, L4977 ); 
   nand2 U1600 ( L4973, L4976, L4978 ); 
   inv U1601 ( L5099, L5105 ); 
   nand2 U1602 ( L5357, L5358, L5359 ); 
   nand2 U1603 ( L5347, L5348, L5362 ); 
   inv U1604 ( L5523, L5529 ); 
   inv U1605 ( L5669, L5675 ); 
   buffer U1606 ( L4389, L5932 ); 
   buffer U1607 ( L2391, L5977 ); 
   buffer U1608 ( L4389, L6052 ); 
   inv U1609 ( L6057, L6063 ); 
   buffer U1610 ( L2635, L6115 ); 
   nor2 U1611 ( L3682, L4389, L6173 ); 
   buffer U1612 ( L3335, L6679 ); 
   inv U1613 ( L6745, L6751 ); 
   inv U1614 ( L6748, L6752 ); 
   inv U1615 ( L6755, L6761 ); 
   inv U1616 ( L6758, L6762 ); 
   inv U1617 ( L6789, L6795 ); 
   inv U1618 ( L6792, L6796 ); 
   inv U1619 ( L6799, L6805 ); 
   inv U1620 ( L6802, L6806 ); 
   inv U1621 ( L6925, L6931 ); 
   buffer U1622 ( L3891, L6983 ); 
   inv U1623 ( L7041, L7047 ); 
   buffer U1624 ( L3979, L7129 ); 
   inv U1625 ( L7273, L7279 ); 
   inv U1626 ( L7276, L7280 ); 
   inv U1627 ( L7283, L7289 ); 
   inv U1628 ( L7286, L7290 ); 
   nand2 U1629 ( L7247, L7248, L7337 ); 
   nand2 U1630 ( L7237, L7238, L7340 ); 
   nand2 U1631 ( L7335, L7336, L7353 ); 
   nand2 U1632 ( L7325, L7326, L7356 ); 
   inv U1633 ( L7531, L7537 ); 
   inv U1634 ( L7534, L7538 ); 
   inv U1635 ( L7541, L7547 ); 
   inv U1636 ( L7544, L7548 ); 
   inv U1637 ( L7575, L7581 ); 
   inv U1638 ( L7578, L7582 ); 
   inv U1639 ( L7585, L7591 ); 
   inv U1640 ( L7588, L7592 ); 
   nand2 U1641 ( L7505, L7506, L7595 ); 
   nand2 U1642 ( L7495, L7496, L7598 ); 
   nand2 U1643 ( L5865, L5872, L2342 ); 
   nand2 U1644 ( L5873, L5880, L2353 ); 
   nand2 U1645 ( L5881, L5888, L2371 ); 
   nand2 U1646 ( L5889, L5896, L2399 ); 
   nand2 U1647 ( L5897, L5904, L2408 ); 
   nand2 U1648 ( L5905, L5912, L2419 ); 
   nand2 U1649 ( L5913, L5920, L2435 ); 
   nand2 U1650 ( L5921, L5928, L2453 ); 
   nand2 U1651 ( L5985, L5992, L2588 ); 
   nand2 U1652 ( L5993, L6000, L2599 ); 
   nand2 U1653 ( L6001, L6008, L2617 ); 
   nand2 U1654 ( L6009, L6016, L2642 ); 
   nand2 U1655 ( L6017, L6024, L2654 ); 
   nand2 U1656 ( L6025, L6032, L2675 ); 
   nand2 U1657 ( L6033, L6040, L2700 ); 
   nand2 U1658 ( L6041, L6048, L2733 ); 
   nand2 U1659 ( L6442, L6445, L3050 ); 
   nand2 U1660 ( L6450, L6453, L3060 ); 
   nand2 U1661 ( L6458, L6461, L3069 ); 
   nand2 U1662 ( L6466, L6469, L3080 ); 
   nand2 U1663 ( L6474, L6477, L3091 ); 
   nand2 U1664 ( L6471, L6478, L3092 ); 
   nand2 U1665 ( L6482, L6485, L3100 ); 
   nand2 U1666 ( L6479, L6486, L3101 ); 
   nand2 U1667 ( L6490, L6493, L3108 ); 
   nand2 U1668 ( L6487, L6494, L3109 ); 
   nand2 U1669 ( L6498, L6501, L3117 ); 
   nand2 U1670 ( L6506, L6509, L3120 ); 
   nand2 U1671 ( L6503, L6510, L3121 ); 
   nand2 U1672 ( L6567, L6574, L3282 ); 
   nand2 U1673 ( L6575, L6582, L3294 ); 
   nand2 U1674 ( L6583, L6590, L3313 ); 
   nand2 U1675 ( L6591, L6598, L3343 ); 
   nand2 U1676 ( L6599, L6606, L3352 ); 
   nand2 U1677 ( L6607, L6614, L3364 ); 
   nand2 U1678 ( L6615, L6622, L3380 ); 
   nand2 U1679 ( L6623, L6630, L3398 ); 
   nand2 U1680 ( L6631, L6638, L3416 ); 
   nand2 U1681 ( L6724, L6727, L3525 ); 
   nand2 U1682 ( L6732, L6735, L3534 ); 
   nand2 U1683 ( L6729, L6736, L3535 ); 
   nand2 U1684 ( L6740, L6743, L3543 ); 
   nand2 U1685 ( L6737, L6744, L3544 ); 
   nand2 U1686 ( L6768, L6771, L3548 ); 
   nand2 U1687 ( L6776, L6779, L3557 ); 
   nand2 U1688 ( L6773, L6780, L3558 ); 
   nand2 U1689 ( L6784, L6787, L3566 ); 
   nand2 U1690 ( L6781, L6788, L3567 ); 
   nand2 U1691 ( L6853, L6860, L3844 ); 
   nand2 U1692 ( L6861, L6868, L3855 ); 
   nand2 U1693 ( L6869, L6876, L3873 ); 
   nand2 U1694 ( L6877, L6884, L3898 ); 
   nand2 U1695 ( L6885, L6892, L3910 ); 
   nand2 U1696 ( L6893, L6900, L3931 ); 
   nand2 U1697 ( L6901, L6908, L3956 ); 
   nand2 U1698 ( L6909, L6916, L3988 ); 
   nand2 U1699 ( L6917, L6924, L3996 ); 
   nand2 U1700 ( L7208, L7211, L4178 ); 
   nand2 U1701 ( L7216, L7219, L4187 ); 
   nand2 U1702 ( L7213, L7220, L4188 ); 
   nand2 U1703 ( L7221, L7228, L4197 ); 
   nand2 U1704 ( L7268, L7271, L4219 ); 
   nand2 U1705 ( L7364, L7367, L4289 ); 
   nand2 U1706 ( L7361, L7368, L4290 ); 
   nand2 U1707 ( L7372, L7375, L4298 ); 
   nand2 U1708 ( L7369, L7376, L4299 ); 
   nand2 U1709 ( L7380, L7383, L4306 ); 
   nand2 U1710 ( L7377, L7384, L4307 ); 
   nand2 U1711 ( L7388, L7391, L4315 ); 
   nand2 U1712 ( L7385, L7392, L4316 ); 
   nand2 U1713 ( L7396, L7399, L4325 ); 
   nand2 U1714 ( L7404, L7407, L4334 ); 
   nand2 U1715 ( L7412, L7415, L4342 ); 
   nand2 U1716 ( L7420, L7423, L4350 ); 
   nand2 U1717 ( L7417, L7424, L4351 ); 
   nand2 U1718 ( L7425, L7432, L4354 ); 
   nand2 U1719 ( L7518, L7521, L4561 ); 
   nand2 U1720 ( L7515, L7522, L4562 ); 
   nand2 U1721 ( L7526, L7529, L4570 ); 
   nand2 U1722 ( L7523, L7530, L4571 ); 
   nand2 U1723 ( L7554, L7557, L4575 ); 
   nand2 U1724 ( L7562, L7565, L4584 ); 
   nand2 U1725 ( L7559, L7566, L4585 ); 
   nand2 U1726 ( L7570, L7573, L4593 ); 
   nand2 U1727 ( L7567, L7574, L4594 ); 
   nand2 U1728 ( L4929, L4936, L4938 ); 
   nand2 U1729 ( L4970, L4977, L4979 ); 
   nand2 U1730 ( L6748, L6751, L6753 ); 
   nand2 U1731 ( L6745, L6752, L6754 ); 
   nand2 U1732 ( L6758, L6761, L6763 ); 
   nand2 U1733 ( L6755, L6762, L6764 ); 
   nand2 U1734 ( L6792, L6795, L6797 ); 
   nand2 U1735 ( L6789, L6796, L6798 ); 
   nand2 U1736 ( L6802, L6805, L6807 ); 
   nand2 U1737 ( L6799, L6806, L6808 ); 
   nand2 U1738 ( L7276, L7279, L7281 ); 
   nand2 U1739 ( L7273, L7280, L7282 ); 
   nand2 U1740 ( L7286, L7289, L7291 ); 
   nand2 U1741 ( L7283, L7290, L7292 ); 
   nand2 U1742 ( L7534, L7537, L7539 ); 
   nand2 U1743 ( L7531, L7538, L7540 ); 
   nand2 U1744 ( L7544, L7547, L7549 ); 
   nand2 U1745 ( L7541, L7548, L7550 ); 
   nand2 U1746 ( L7578, L7581, L7583 ); 
   nand2 U1747 ( L7575, L7582, L7584 ); 
   nand2 U1748 ( L7588, L7591, L7593 ); 
   nand2 U1749 ( L7585, L7592, L7594 ); 
   inv U1750 ( L1850, L1856 ); 
   and5 U1751 ( L895, L853, L827, L805, L792, L920 ); 
   and2 U1752 ( L792, L821, L925 ); 
   and3 U1753 ( L805, L792, L845, L926 ); 
   and4 U1754 ( L827, L792, L868, L805, L927 ); 
   and5 U1755 ( L853, L827, L792, L877, L805, L928 ); 
   and2 U1756 ( L805, L845, L937 ); 
   and3 U1757 ( L827, L868, L805, L938 ); 
   and4 U1758 ( L853, L827, L877, L805, L939 ); 
   and4 U1759 ( L895, L827, L805, L853, L940 ); 
   and2 U1760 ( L805, L845, L941 ); 
   and3 U1761 ( L827, L868, L805, L942 ); 
   and4 U1762 ( L853, L827, L877, L805, L943 ); 
   and2 U1763 ( L827, L868, L944 ); 
   and3 U1764 ( L853, L827, L877, L945 ); 
   and3 U1765 ( L895, L827, L853, L946 ); 
   and2 U1766 ( L827, L868, L947 ); 
   and3 U1767 ( L853, L827, L877, L948 ); 
   and2 U1768 ( L853, L877, L949 ); 
   and2 U1769 ( L895, L853, L956 ); 
   and5 U1770 ( L1038, L1093, L1055, L1026, L1074, L1122 ); 
   and2 U1771 ( L1026, L1050, L1125 ); 
   and3 U1772 ( L1038, L1026, L1068, L1126 ); 
   and4 U1773 ( L1055, L1026, L1086, L1038, L1127 ); 
   and5 U1774 ( L1074, L1055, L1026, L1102, L1038, L1128 ); 
   and2 U1775 ( L1038, L1068, L1132 ); 
   and3 U1776 ( L1055, L1086, L1038, L1133 ); 
   and4 U1777 ( L1074, L1055, L1102, L1038, L1134 ); 
   and2 U1778 ( L1086, L1055, L1137 ); 
   and3 U1779 ( L1074, L1055, L1102, L1138 ); 
   and2 U1780 ( L1074, L1102, L1141 ); 
   inv U1781 ( L1217, L1221 ); 
   inv U1782 ( L1226, L1230 ); 
   inv U1783 ( L1240, L1244 ); 
   inv U1784 ( L1249, L1253 ); 
   inv U1785 ( L1263, L1267 ); 
   inv U1786 ( L1272, L1276 ); 
   buffer U1787 ( L1235, L1284 ); 
   buffer U1788 ( L1235, L1288 ); 
   buffer U1789 ( L1258, L1292 ); 
   buffer U1790 ( L1258, L1296 ); 
   buffer U1791 ( L1281, L1300 ); 
   buffer U1792 ( L1281, L1304 ); 
   and4 U1793 ( L1687, L1573, L1556, L1546, L1702 ); 
   and2 U1794 ( L1546, L1567, L1705 ); 
   and3 U1795 ( L1556, L1546, L1584, L1706 ); 
   and4 U1796 ( L1573, L1546, L1590, L1556, L1707 ); 
   and2 U1797 ( L1556, L1584, L1709 ); 
   and3 U1798 ( L1573, L1590, L1556, L1710 ); 
   and3 U1799 ( L1687, L1573, L1556, L1711 ); 
   and2 U1800 ( L1556, L1584, L1712 ); 
   and3 U1801 ( L1573, L1590, L1556, L1713 ); 
   and2 U1802 ( L1573, L1590, L1714 ); 
   and5 U1803 ( L1695, L1655, L1630, L1609, L1598, L1718 ); 
   and2 U1804 ( L1598, L1624, L1722 ); 
   and3 U1805 ( L1609, L1598, L1647, L1723 ); 
   and4 U1806 ( L1630, L1598, L1669, L1609, L1724 ); 
   and5 U1807 ( L1655, L1630, L1598, L1677, L1609, L1725 ); 
   and2 U1808 ( L1609, L1647, L1733 ); 
   and3 U1809 ( L1630, L1669, L1609, L1734 ); 
   and4 U1810 ( L1655, L1630, L1677, L1609, L1735 ); 
   and4 U1811 ( L1695, L1630, L1609, L1655, L1736 ); 
   and2 U1812 ( L1609, L1647, L1737 ); 
   and3 U1813 ( L1630, L1669, L1609, L1738 ); 
   and4 U1814 ( L1655, L1630, L1677, L1609, L1739 ); 
   and2 U1815 ( L1630, L1669, L1740 ); 
   and3 U1816 ( L1655, L1630, L1677, L1741 ); 
   and3 U1817 ( L1695, L1630, L1655, L1742 ); 
   and2 U1818 ( L1630, L1669, L1743 ); 
   and3 U1819 ( L1655, L1630, L1677, L1744 ); 
   and2 U1820 ( L1655, L1677, L1745 ); 
   and2 U1821 ( L1687, L1573, L1749 ); 
   and2 U1822 ( L1695, L1655, L1750 ); 
   and4 U1823 ( L1805, L1850, L1822, L1795, L1935 ); 
   and2 U1824 ( L1795, L1816, L1938 ); 
   and3 U1825 ( L1805, L1795, L1834, L1939 ); 
   and4 U1826 ( L1822, L1795, L1841, L1805, L1940 ); 
   and2 U1827 ( L1805, L1834, L1942 ); 
   and3 U1828 ( L1822, L1841, L1805, L1943 ); 
   and3 U1829 ( L1850, L1822, L1805, L1944 ); 
   and2 U1830 ( L1805, L1834, L1945 ); 
   and3 U1831 ( L1841, L1822, L1805, L1946 ); 
   and2 U1832 ( L1822, L1841, L1947 ); 
   and2 U1833 ( L1850, L1822, L1948 ); 
   and2 U1834 ( L1822, L1841, L1949 ); 
   and5 U1835 ( L1869, L1921, L1885, L1859, L1903, L1950 ); 
   and2 U1836 ( L1859, L1880, L1953 ); 
   and3 U1837 ( L1869, L1859, L1897, L1954 ); 
   and4 U1838 ( L1885, L1859, L1914, L1869, L1955 ); 
   and5 U1839 ( L1903, L1885, L1859, L1929, L1869, L1956 ); 
   and2 U1840 ( L1869, L1897, L1960 ); 
   and3 U1841 ( L1885, L1914, L1869, L1961 ); 
   and4 U1842 ( L1903, L1885, L1929, L1869, L1962 ); 
   and2 U1843 ( L1914, L1885, L1965 ); 
   and3 U1844 ( L1903, L1885, L1929, L1966 ); 
   and2 U1845 ( L1903, L1929, L1969 ); 
   nand2 U1846 ( L2341, L2342, L2343 ); 
   nand2 U1847 ( L2352, L2353, L2354 ); 
   nand2 U1848 ( L2370, L2371, L2372 ); 
   nand2 U1849 ( L2398, L2399, L2400 ); 
   nand2 U1850 ( L2407, L2408, L2409 ); 
   nand2 U1851 ( L2418, L2419, L2420 ); 
   nand2 U1852 ( L2434, L2435, L2436 ); 
   nand2 U1853 ( L2452, L2453, L2454 ); 
   nand2 U1854 ( L5932, L5935, L2470 ); 
   inv U1855 ( L5932, L5936 ); 
   inv U1856 ( L5977, L5983 ); 
   nand2 U1857 ( L2587, L2588, L2589 ); 
   nand2 U1858 ( L2598, L2599, L2600 ); 
   nand2 U1859 ( L2616, L2617, L2618 ); 
   nand2 U1860 ( L2641, L2642, L2643 ); 
   nand2 U1861 ( L2653, L2654, L2655 ); 
   nand2 U1862 ( L2674, L2675, L2676 ); 
   nand2 U1863 ( L2699, L2700, L2701 ); 
   nand2 U1864 ( L2732, L2733, L2734 ); 
   nand2 U1865 ( L6052, L6055, L2740 ); 
   inv U1866 ( L6052, L6056 ); 
   and4 U1867 ( L3018, L2973, L2965, L2956, L3022 ); 
   and2 U1868 ( L2956, L2970, L3025 ); 
   and3 U1869 ( L2965, L2956, L2977, L3026 ); 
   and4 U1870 ( L2973, L2956, L2979, L2965, L3027 ); 
   and5 U1871 ( L3021, L3009, L3001, L2992, L2982, L3029 ); 
   and2 U1872 ( L2982, L2998, L3030 ); 
   and3 U1873 ( L2992, L2982, L3006, L3031 ); 
   and4 U1874 ( L3001, L2982, L3013, L2992, L3032 ); 
   and5 U1875 ( L3009, L3001, L2982, L3015, L2992, L3033 ); 
   nand2 U1876 ( L3050, L3051, L3052 ); 
   nand2 U1877 ( L3060, L3061, L3062 ); 
   nand2 U1878 ( L3069, L3070, L3071 ); 
   nand2 U1879 ( L3080, L3081, L3082 ); 
   nand2 U1880 ( L3091, L3092, L3093 ); 
   nand2 U1881 ( L3100, L3101, L3102 ); 
   nand2 U1882 ( L3108, L3109, L3110 ); 
   nand2 U1883 ( L3117, L3118, L3119 ); 
   nand2 U1884 ( L3120, L3121, L3122 ); 
   and5 U1885 ( L3215, L3203, L3195, L3186, L3176, L3228 ); 
   and2 U1886 ( L3176, L3192, L3231 ); 
   and3 U1887 ( L3186, L3176, L3200, L3232 ); 
   and4 U1888 ( L3195, L3176, L3207, L3186, L3233 ); 
   and5 U1889 ( L3203, L3195, L3176, L3209, L3186, L3234 ); 
   nand2 U1890 ( L3281, L3282, L3283 ); 
   nand2 U1891 ( L3293, L3294, L3295 ); 
   nand2 U1892 ( L3312, L3313, L3314 ); 
   nand2 U1893 ( L3342, L3343, L3344 ); 
   nand2 U1894 ( L3351, L3352, L3353 ); 
   nand2 U1895 ( L3363, L3364, L3365 ); 
   nand2 U1896 ( L3379, L3380, L3381 ); 
   nand2 U1897 ( L3397, L3398, L3399 ); 
   nand2 U1898 ( L3415, L3416, L3417 ); 
   inv U1899 ( L6679, L6685 ); 
   inv U1900 ( L3504, L3508 ); 
   inv U1901 ( L3513, L3517 ); 
   nand2 U1902 ( L3525, L3526, L3527 ); 
   nand2 U1903 ( L3534, L3535, L3536 ); 
   nand2 U1904 ( L3543, L3544, L3545 ); 
   nand2 U1905 ( L3548, L3549, L3550 ); 
   nand2 U1906 ( L3557, L3558, L3559 ); 
   nand2 U1907 ( L3566, L3567, L3568 ); 
   buffer U1908 ( L3522, L3571 ); 
   buffer U1909 ( L3522, L3575 ); 
   nand2 U1910 ( L3843, L3844, L3845 ); 
   nand2 U1911 ( L3854, L3855, L3856 ); 
   nand2 U1912 ( L3872, L3873, L3874 ); 
   nand2 U1913 ( L3897, L3898, L3899 ); 
   nand2 U1914 ( L3909, L3910, L3911 ); 
   nand2 U1915 ( L3930, L3931, L3932 ); 
   nand2 U1916 ( L3955, L3956, L3957 ); 
   nand2 U1917 ( L3987, L3988, L3989 ); 
   nand2 U1918 ( L3995, L3996, L3997 ); 
   nand2 U1919 ( L4178, L4179, L4180 ); 
   nand2 U1920 ( L4187, L4188, L4189 ); 
   nand2 U1921 ( L4196, L4197, L4198 ); 
   inv U1922 ( L4203, L4207 ); 
   inv U1923 ( L4212, L4216 ); 
   nand2 U1924 ( L4219, L4220, L4221 ); 
   inv U1925 ( L4226, L4230 ); 
   inv U1926 ( L4235, L4239 ); 
   buffer U1927 ( L4244, L4263 ); 
   buffer U1928 ( L4244, L4267 ); 
   nand2 U1929 ( L4289, L4290, L4291 ); 
   nand2 U1930 ( L4298, L4299, L4300 ); 
   nand2 U1931 ( L4306, L4307, L4308 ); 
   nand2 U1932 ( L4315, L4316, L4317 ); 
   nand2 U1933 ( L4325, L4326, L4327 ); 
   nand2 U1934 ( L4334, L4335, L4336 ); 
   nand2 U1935 ( L4342, L4343, L4344 ); 
   nand2 U1936 ( L4350, L4351, L4352 ); 
   nand2 U1937 ( L4353, L4354, L4355 ); 
   inv U1938 ( L4531, L4535 ); 
   inv U1939 ( L4540, L4544 ); 
   inv U1940 ( L4554, L4558 ); 
   nand2 U1941 ( L4561, L4562, L4563 ); 
   nand2 U1942 ( L4570, L4571, L4572 ); 
   nand2 U1943 ( L4575, L4576, L4577 ); 
   nand2 U1944 ( L4584, L4585, L4586 ); 
   nand2 U1945 ( L4593, L4594, L4595 ); 
   buffer U1946 ( L4549, L4598 ); 
   buffer U1947 ( L4549, L4602 ); 
   buffer U1948 ( L1921, L4716 ); 
   buffer U1949 ( L1859, L4724 ); 
   buffer U1950 ( L1869, L4732 ); 
   buffer U1951 ( L1885, L4740 ); 
   buffer U1952 ( L1903, L4748 ); 
   buffer U1953 ( L1093, L4756 ); 
   buffer U1954 ( L1026, L4764 ); 
   buffer U1955 ( L1038, L4772 ); 
   buffer U1956 ( L1055, L4780 ); 
   buffer U1957 ( L1074, L4788 ); 
   nand2 U1958 ( L4937, L4938, L4939 ); 
   nand2 U1959 ( L4978, L4979, L4980 ); 
   buffer U1960 ( L895, L5044 ); 
   buffer U1961 ( L853, L5054 ); 
   buffer U1962 ( L792, L5064 ); 
   buffer U1963 ( L827, L5074 ); 
   buffer U1964 ( L805, L5084 ); 
   buffer U1965 ( L805, L5094 ); 
   buffer U1966 ( L895, L5132 ); 
   buffer U1967 ( L853, L5142 ); 
   buffer U1968 ( L792, L5152 ); 
   buffer U1969 ( L827, L5162 ); 
   inv U1970 ( L5359, L5365 ); 
   inv U1971 ( L5362, L5366 ); 
   buffer U1972 ( L1687, L5488 ); 
   buffer U1973 ( L1573, L5498 ); 
   buffer U1974 ( L1546, L5508 ); 
   buffer U1975 ( L1556, L5518 ); 
   buffer U1976 ( L1687, L5546 ); 
   buffer U1977 ( L1573, L5556 ); 
   buffer U1978 ( L1546, L5566 ); 
   buffer U1979 ( L1556, L5576 ); 
   buffer U1980 ( L1695, L5614 ); 
   buffer U1981 ( L1655, L5624 ); 
   buffer U1982 ( L1598, L5634 ); 
   buffer U1983 ( L1630, L5644 ); 
   buffer U1984 ( L1609, L5654 ); 
   buffer U1985 ( L1609, L5664 ); 
   buffer U1986 ( L1695, L5702 ); 
   buffer U1987 ( L1655, L5712 ); 
   buffer U1988 ( L1598, L5722 ); 
   buffer U1989 ( L1630, L5732 ); 
   buffer U1990 ( L1795, L5820 ); 
   buffer U1991 ( L1795, L5828 ); 
   buffer U1992 ( L1805, L5836 ); 
   buffer U1993 ( L1805, L5844 ); 
   buffer U1994 ( L1822, L5852 ); 
   buffer U1995 ( L1822, L5860 ); 
   inv U1996 ( L6115, L6121 ); 
   inv U1997 ( L6173, L6179 ); 
   buffer U1998 ( L2724, L6261 ); 
   inv U1999 ( L7353, L7359 ); 
   inv U2000 ( L7356, L7360 ); 
   inv U2001 ( L7337, L7343 ); 
   inv U2002 ( L7340, L7344 ); 
   nand2 U2003 ( L6763, L6764, L6809 ); 
   nand2 U2004 ( L6753, L6754, L6812 ); 
   nand2 U2005 ( L6807, L6808, L6819 ); 
   nand2 U2006 ( L6797, L6798, L6822 ); 
   inv U2007 ( L6983, L6989 ); 
   inv U2008 ( L7129, L7135 ); 
   nand2 U2009 ( L7291, L7292, L7345 ); 
   nand2 U2010 ( L7281, L7282, L7348 ); 
   inv U2011 ( L7595, L7601 ); 
   inv U2012 ( L7598, L7602 ); 
   nand2 U2013 ( L7549, L7550, L7603 ); 
   nand2 U2014 ( L7539, L7540, L7606 ); 
   nand2 U2015 ( L7593, L7594, L7611 ); 
   nand2 U2016 ( L7583, L7584, L7614 ); 
   or5 U2017 ( L802, L925, L926, L927, L928, L929 ); 
   or2 U2018 ( L868, L949, L950 ); 
   or5 U2019 ( L1035, L1125, L1126, L1127, L1128, L1129 ); 
   or4 U2020 ( L1553, L1705, L1706, L1707, L1708 ); 
   or2 U2021 ( L1584, L1714, L1715 ); 
   or5 U2022 ( L1606, L1722, L1723, L1724, L1725, L1726 ); 
   or2 U2023 ( L1669, L1745, L1746 ); 
   or4 U2024 ( L1802, L1938, L1939, L1940, L1941 ); 
   or5 U2025 ( L1866, L1953, L1954, L1955, L1956, L1957 ); 
   nand2 U2026 ( L5929, L5936, L2471 ); 
   nand2 U2027 ( L6049, L6056, L2741 ); 
   or4 U2028 ( L2962, L3025, L3026, L3027, L3028 ); 
   or5 U2029 ( L2989, L3030, L3031, L3032, L3033, L3034 ); 
   or5 U2030 ( L3183, L3231, L3232, L3233, L3234, L3235 ); 
   or4 U2031 ( L845, L944, L945, L946, L5014 ); 
   or5 U2032 ( L821, L937, L938, L939, L940, L5034 ); 
   nor3 U2033 ( L845, L947, L948, L5102 ); 
   nor4 U2034 ( L821, L941, L942, L943, L5122 ); 
   nand2 U2035 ( L5362, L5365, L5367 ); 
   nand2 U2036 ( L5359, L5366, L5368 ); 
   or4 U2037 ( L1567, L1709, L1710, L1711, L5478 ); 
   nor3 U2038 ( L1567, L1712, L1713, L5536 ); 
   or4 U2039 ( L1647, L1740, L1741, L1742, L5584 ); 
   or5 U2040 ( L1624, L1733, L1734, L1735, L1736, L5604 ); 
   nor3 U2041 ( L1647, L1743, L1744, L5672 ); 
   nor4 U2042 ( L1624, L1737, L1738, L1739, L5692 ); 
   or4 U2043 ( L1816, L1942, L1943, L1944, L5817 ); 
   nor3 U2044 ( L1816, L1945, L1946, L5825 ); 
   or3 U2045 ( L1834, L1947, L1948, L5833 ); 
   nor2 U2046 ( L1834, L1949, L5841 ); 
   nand2 U2047 ( L7356, L7359, L6340 ); 
   nand2 U2048 ( L7353, L7360, L6341 ); 
   nand2 U2049 ( L7340, L7343, L6350 ); 
   nand2 U2050 ( L7337, L7344, L6351 ); 
   nand2 U2051 ( L7598, L7601, L7436 ); 
   nand2 U2052 ( L7595, L7602, L7437 ); 
   inv U2053 ( L4716, L4720 ); 
   inv U2054 ( L4724, L4728 ); 
   inv U2055 ( L4732, L4736 ); 
   inv U2056 ( L4740, L4744 ); 
   inv U2057 ( L4748, L4752 ); 
   inv U2058 ( L4756, L4760 ); 
   inv U2059 ( L4764, L4768 ); 
   inv U2060 ( L4772, L4776 ); 
   inv U2061 ( L4780, L4784 ); 
   inv U2062 ( L4788, L4792 ); 
   inv U2063 ( L3344, L3350 ); 
   inv U2064 ( L2400, L2406 ); 
   inv U2065 ( L920, L924 ); 
   inv U2066 ( L5084, L5088 ); 
   inv U2067 ( L5094, L5098 ); 
   and2 U2068 ( L902, L920, L997 ); 
   and2 U2069 ( L1108, L1122, L1146 ); 
   inv U2070 ( L1284, L1287 ); 
   inv U2071 ( L1288, L1291 ); 
   inv U2072 ( L1292, L1295 ); 
   inv U2073 ( L1296, L1299 ); 
   inv U2074 ( L1300, L1303 ); 
   inv U2075 ( L1304, L1307 ); 
   and3 U2076 ( L1226, L1217, L1284, L1309 ); 
   and3 U2077 ( L1230, L1221, L1288, L1312 ); 
   and3 U2078 ( L1249, L1240, L1292, L1315 ); 
   and3 U2079 ( L1253, L1244, L1296, L1318 ); 
   and3 U2080 ( L1272, L1263, L1300, L1321 ); 
   and3 U2081 ( L1276, L1267, L1304, L1324 ); 
   inv U2082 ( L1718, L1721 ); 
   inv U2083 ( L5518, L5522 ); 
   inv U2084 ( L5576, L5580 ); 
   inv U2085 ( L5654, L5658 ); 
   inv U2086 ( L5664, L5668 ); 
   and2 U2087 ( L1702, L1718, L1788 ); 
   and2 U2088 ( L1935, L1950, L1974 ); 
   inv U2089 ( L5820, L5824 ); 
   inv U2090 ( L5828, L5832 ); 
   inv U2091 ( L5836, L5840 ); 
   inv U2092 ( L5844, L5848 ); 
   nand2 U2093 ( L5852, L5855, L1999 ); 
   inv U2094 ( L5852, L5856 ); 
   nand2 U2095 ( L5860, L5863, L2003 ); 
   inv U2096 ( L5860, L5864 ); 
   nand2 U2097 ( L2470, L2471, L2472 ); 
   and4 U2098 ( L2354, L2400, L2372, L2343, L2487 ); 
   and2 U2099 ( L2343, L2366, L2492 ); 
   and3 U2100 ( L2354, L2343, L2384, L2493 ); 
   and4 U2101 ( L2372, L2343, L2391, L2354, L2494 ); 
   and2 U2102 ( L2354, L2384, L2500 ); 
   and3 U2103 ( L2372, L2391, L2354, L2501 ); 
   and3 U2104 ( L2400, L2372, L2354, L2502 ); 
   and2 U2105 ( L2354, L2384, L2503 ); 
   and3 U2106 ( L2391, L2372, L2354, L2504 ); 
   and2 U2107 ( L2372, L2391, L2505 ); 
   and2 U2108 ( L2400, L2372, L2506 ); 
   and2 U2109 ( L2372, L2391, L2507 ); 
   and2 U2110 ( L2409, L2431, L2511 ); 
   and3 U2111 ( L2420, L2409, L2448, L2512 ); 
   and4 U2112 ( L2436, L2409, L2465, L2420, L2513 ); 
   and5 U2113 ( L2454, L2436, L2409, L2481, L2420, L2514 ); 
   and2 U2114 ( L2420, L2448, L2518 ); 
   and3 U2115 ( L2436, L2465, L2420, L2519 ); 
   and4 U2116 ( L2454, L2436, L2481, L2420, L2520 ); 
   and2 U2117 ( L2465, L2436, L2523 ); 
   and3 U2118 ( L2454, L2436, L2481, L2524 ); 
   and2 U2119 ( L2454, L2481, L2527 ); 
   nand2 U2120 ( L2740, L2741, L2742 ); 
   and4 U2121 ( L2734, L2618, L2600, L2589, L2749 ); 
   and2 U2122 ( L2589, L2612, L2754 ); 
   and3 U2123 ( L2600, L2589, L2629, L2755 ); 
   and4 U2124 ( L2618, L2589, L2635, L2600, L2756 ); 
   and2 U2125 ( L2600, L2629, L2762 ); 
   and3 U2126 ( L2618, L2635, L2600, L2763 ); 
   and3 U2127 ( L2734, L2618, L2600, L2764 ); 
   and2 U2128 ( L2600, L2629, L2765 ); 
   and3 U2129 ( L2618, L2635, L2600, L2766 ); 
   and2 U2130 ( L2618, L2635, L2767 ); 
   and2 U2131 ( L2643, L2670, L2776 ); 
   and3 U2132 ( L2655, L2643, L2693, L2777 ); 
   and4 U2133 ( L2676, L2643, L2715, L2655, L2778 ); 
   and5 U2134 ( L2701, L2676, L2643, L2724, L2655, L2779 ); 
   and2 U2135 ( L2655, L2693, L2788 ); 
   and3 U2136 ( L2676, L2715, L2655, L2789 ); 
   and4 U2137 ( L2701, L2676, L2724, L2655, L2790 ); 
   and2 U2138 ( L2655, L2693, L2792 ); 
   and3 U2139 ( L2676, L2715, L2655, L2793 ); 
   and4 U2140 ( L2701, L2676, L2724, L2655, L2794 ); 
   and2 U2141 ( L2676, L2715, L2795 ); 
   and3 U2142 ( L2701, L2676, L2724, L2796 ); 
   and2 U2143 ( L2676, L2715, L2798 ); 
   and3 U2144 ( L2701, L2676, L2724, L2799 ); 
   and2 U2145 ( L2701, L2724, L2800 ); 
   and2 U2146 ( L2734, L2618, L2804 ); 
   and2 U2147 ( L3022, L3029, L3035 ); 
   and2 U2148 ( L3022, L3034, L3045 ); 
   and4 U2149 ( L3119, L3071, L3062, L3052, L3123 ); 
   and2 U2150 ( L3052, L3068, L3128 ); 
   and3 U2151 ( L3062, L3052, L3076, L3129 ); 
   and4 U2152 ( L3071, L3052, L3079, L3062, L3130 ); 
   and5 U2153 ( L3122, L3110, L3102, L3093, L3082, L3136 ); 
   and2 U2154 ( L3082, L3099, L3139 ); 
   and3 U2155 ( L3093, L3082, L3107, L3140 ); 
   and4 U2156 ( L3102, L3082, L3114, L3093, L3141 ); 
   and5 U2157 ( L3110, L3102, L3082, L3116, L3093, L3142 ); 
   and2 U2158 ( L3216, L3228, L3249 ); 
   and4 U2159 ( L3295, L3344, L3314, L3283, L3431 ); 
   and2 U2160 ( L3283, L3308, L3434 ); 
   and3 U2161 ( L3295, L3283, L3327, L3435 ); 
   and4 U2162 ( L3314, L3283, L3335, L3295, L3436 ); 
   and2 U2163 ( L3295, L3327, L3438 ); 
   and3 U2164 ( L3314, L3335, L3295, L3439 ); 
   and3 U2165 ( L3344, L3314, L3295, L3440 ); 
   and2 U2166 ( L3295, L3327, L3441 ); 
   and3 U2167 ( L3335, L3314, L3295, L3442 ); 
   and2 U2168 ( L3314, L3335, L3443 ); 
   and2 U2169 ( L3344, L3314, L3444 ); 
   and2 U2170 ( L3314, L3335, L3445 ); 
   and5 U2171 ( L3365, L3417, L3381, L3353, L3399, L3446 ); 
   and2 U2172 ( L3353, L3376, L3449 ); 
   and3 U2173 ( L3365, L3353, L3393, L3450 ); 
   and4 U2174 ( L3381, L3353, L3410, L3365, L3451 ); 
   and5 U2175 ( L3399, L3381, L3353, L3425, L3365, L3452 ); 
   and2 U2176 ( L3365, L3393, L3456 ); 
   and3 U2177 ( L3381, L3410, L3365, L3457 ); 
   and4 U2178 ( L3399, L3381, L3425, L3365, L3458 ); 
   and2 U2179 ( L3410, L3381, L3460 ); 
   and3 U2180 ( L3399, L3381, L3425, L3461 ); 
   and2 U2181 ( L3399, L3425, L3463 ); 
   inv U2182 ( L3527, L3531 ); 
   inv U2183 ( L3536, L3540 ); 
   inv U2184 ( L3550, L3554 ); 
   inv U2185 ( L3559, L3563 ); 
   inv U2186 ( L3571, L3574 ); 
   inv U2187 ( L3575, L3578 ); 
   buffer U2188 ( L3545, L3579 ); 
   buffer U2189 ( L3545, L3583 ); 
   buffer U2190 ( L3568, L3587 ); 
   buffer U2191 ( L3568, L3591 ); 
   and3 U2192 ( L3513, L3504, L3571, L3596 ); 
   and3 U2193 ( L3517, L3508, L3575, L3599 ); 
   and4 U2194 ( L3989, L3874, L3856, L3845, L4004 ); 
   and2 U2195 ( L3845, L3868, L4007 ); 
   and3 U2196 ( L3856, L3845, L3885, L4008 ); 
   and4 U2197 ( L3874, L3845, L3891, L3856, L4009 ); 
   and2 U2198 ( L3856, L3885, L4011 ); 
   and3 U2199 ( L3874, L3891, L3856, L4012 ); 
   and3 U2200 ( L3989, L3874, L3856, L4013 ); 
   and2 U2201 ( L3856, L3885, L4014 ); 
   and3 U2202 ( L3874, L3891, L3856, L4015 ); 
   and2 U2203 ( L3874, L3891, L4016 ); 
   and5 U2204 ( L3997, L3957, L3932, L3911, L3899, L4020 ); 
   and2 U2205 ( L3899, L3926, L4024 ); 
   and3 U2206 ( L3911, L3899, L3949, L4025 ); 
   and4 U2207 ( L3932, L3899, L3971, L3911, L4026 ); 
   and5 U2208 ( L3957, L3932, L3899, L3979, L3911, L4027 ); 
   and2 U2209 ( L3911, L3949, L4035 ); 
   and3 U2210 ( L3932, L3971, L3911, L4036 ); 
   and4 U2211 ( L3957, L3932, L3979, L3911, L4037 ); 
   and4 U2212 ( L3997, L3932, L3911, L3957, L4038 ); 
   and2 U2213 ( L3911, L3949, L4039 ); 
   and3 U2214 ( L3932, L3971, L3911, L4040 ); 
   and4 U2215 ( L3957, L3932, L3979, L3911, L4041 ); 
   and2 U2216 ( L3932, L3971, L4042 ); 
   and3 U2217 ( L3957, L3932, L3979, L4043 ); 
   and3 U2218 ( L3997, L3932, L3957, L4044 ); 
   and2 U2219 ( L3932, L3971, L4045 ); 
   and3 U2220 ( L3957, L3932, L3979, L4046 ); 
   and2 U2221 ( L3957, L3979, L4047 ); 
   and2 U2222 ( L3989, L3874, L4051 ); 
   and2 U2223 ( L3997, L3957, L4052 ); 
   inv U2224 ( L4180, L4184 ); 
   inv U2225 ( L4189, L4193 ); 
   buffer U2226 ( L4198, L4247 ); 
   buffer U2227 ( L4198, L4251 ); 
   buffer U2228 ( L4221, L4255 ); 
   buffer U2229 ( L4221, L4259 ); 
   inv U2230 ( L4263, L4266 ); 
   inv U2231 ( L4267, L4270 ); 
   and3 U2232 ( L4235, L4226, L4263, L4284 ); 
   and3 U2233 ( L4239, L4230, L4267, L4287 ); 
   and4 U2234 ( L4352, L4308, L4300, L4291, L4356 ); 
   and2 U2235 ( L4291, L4305, L4361 ); 
   and3 U2236 ( L4300, L4291, L4312, L4362 ); 
   and4 U2237 ( L4308, L4291, L4314, L4300, L4363 ); 
   and5 U2238 ( L4355, L4344, L4336, L4327, L4317, L4369 ); 
   and2 U2239 ( L4317, L4333, L4372 ); 
   and3 U2240 ( L4327, L4317, L4341, L4373 ); 
   and4 U2241 ( L4336, L4317, L4348, L4327, L4374 ); 
   and5 U2242 ( L4344, L4336, L4317, L4349, L4327, L4375 ); 
   inv U2243 ( L4563, L4567 ); 
   inv U2244 ( L4577, L4581 ); 
   inv U2245 ( L4586, L4590 ); 
   inv U2246 ( L4598, L4601 ); 
   inv U2247 ( L4602, L4605 ); 
   buffer U2248 ( L4572, L4606 ); 
   buffer U2249 ( L4572, L4610 ); 
   buffer U2250 ( L4595, L4614 ); 
   buffer U2251 ( L4595, L4618 ); 
   and3 U2252 ( L4540, L4531, L4598, L4623 ); 
   and3 U2253 ( L4544, L4535, L4602, L4626 ); 
   buffer U2254 ( L3417, L4796 ); 
   buffer U2255 ( L3353, L4804 ); 
   buffer U2256 ( L3365, L4812 ); 
   buffer U2257 ( L3381, L4820 ); 
   buffer U2258 ( L3399, L4828 ); 
   buffer U2259 ( L2409, L4844 ); 
   buffer U2260 ( L2420, L4852 ); 
   buffer U2261 ( L2436, L4860 ); 
   buffer U2262 ( L2454, L4868 ); 
   inv U2263 ( L4939, L4945 ); 
   nand2 U2264 ( L4939, L4946, L4948 ); 
   inv U2265 ( L4980, L4986 ); 
   nand2 U2266 ( L4980, L4987, L4989 ); 
   inv U2267 ( L5044, L5048 ); 
   inv U2268 ( L5054, L5058 ); 
   inv U2269 ( L5064, L5068 ); 
   inv U2270 ( L5074, L5078 ); 
   inv U2271 ( L5162, L5166 ); 
   inv U2272 ( L5132, L5136 ); 
   inv U2273 ( L5142, L5146 ); 
   inv U2274 ( L5152, L5156 ); 
   nand2 U2275 ( L5367, L5368, L5388 ); 
   inv U2276 ( L5488, L5492 ); 
   inv U2277 ( L5498, L5502 ); 
   inv U2278 ( L5508, L5512 ); 
   inv U2279 ( L5546, L5550 ); 
   inv U2280 ( L5556, L5560 ); 
   inv U2281 ( L5566, L5570 ); 
   inv U2282 ( L5614, L5618 ); 
   inv U2283 ( L5624, L5628 ); 
   inv U2284 ( L5634, L5638 ); 
   inv U2285 ( L5644, L5648 ); 
   inv U2286 ( L5732, L5736 ); 
   inv U2287 ( L5702, L5706 ); 
   inv U2288 ( L5712, L5716 ); 
   inv U2289 ( L5722, L5726 ); 
   buffer U2290 ( L2343, L5940 ); 
   buffer U2291 ( L2343, L5948 ); 
   buffer U2292 ( L2354, L5956 ); 
   buffer U2293 ( L2354, L5964 ); 
   buffer U2294 ( L2372, L5972 ); 
   buffer U2295 ( L2372, L5980 ); 
   buffer U2296 ( L2734, L6080 ); 
   buffer U2297 ( L2618, L6090 ); 
   buffer U2298 ( L2589, L6100 ); 
   buffer U2299 ( L2600, L6110 ); 
   buffer U2300 ( L2734, L6138 ); 
   buffer U2301 ( L2618, L6148 ); 
   buffer U2302 ( L2589, L6158 ); 
   buffer U2303 ( L2600, L6168 ); 
   buffer U2304 ( L2701, L6216 ); 
   buffer U2305 ( L2643, L6226 ); 
   buffer U2306 ( L2676, L6236 ); 
   buffer U2307 ( L2655, L6246 ); 
   buffer U2308 ( L2655, L6256 ); 
   inv U2309 ( L6261, L6267 ); 
   buffer U2310 ( L2701, L6304 ); 
   buffer U2311 ( L2643, L6314 ); 
   buffer U2312 ( L2676, L6324 ); 
   nand2 U2313 ( L6340, L6341, L6342 ); 
   nand2 U2314 ( L6350, L6351, L6352 ); 
   inv U2315 ( L7345, L7351 ); 
   inv U2316 ( L7348, L7352 ); 
   buffer U2317 ( L3283, L6642 ); 
   buffer U2318 ( L3283, L6650 ); 
   buffer U2319 ( L3295, L6658 ); 
   buffer U2320 ( L3295, L6666 ); 
   buffer U2321 ( L3314, L6674 ); 
   buffer U2322 ( L3314, L6682 ); 
   inv U2323 ( L6809, L6815 ); 
   inv U2324 ( L6812, L6816 ); 
   inv U2325 ( L6819, L6825 ); 
   inv U2326 ( L6822, L6826 ); 
   buffer U2327 ( L3989, L6948 ); 
   buffer U2328 ( L3874, L6958 ); 
   buffer U2329 ( L3845, L6968 ); 
   buffer U2330 ( L3856, L6978 ); 
   buffer U2331 ( L3989, L7006 ); 
   buffer U2332 ( L3874, L7016 ); 
   buffer U2333 ( L3845, L7026 ); 
   buffer U2334 ( L3856, L7036 ); 
   buffer U2335 ( L3997, L7074 ); 
   buffer U2336 ( L3957, L7084 ); 
   buffer U2337 ( L3899, L7094 ); 
   buffer U2338 ( L3932, L7104 ); 
   buffer U2339 ( L3911, L7114 ); 
   buffer U2340 ( L3911, L7124 ); 
   buffer U2341 ( L3997, L7162 ); 
   buffer U2342 ( L3957, L7172 ); 
   buffer U2343 ( L3899, L7182 ); 
   buffer U2344 ( L3932, L7192 ); 
   nand2 U2345 ( L7436, L7437, L7438 ); 
   inv U2346 ( L7611, L7617 ); 
   inv U2347 ( L7614, L7618 ); 
   inv U2348 ( L7603, L7609 ); 
   inv U2349 ( L7606, L7610 ); 
   and2 U2350 ( L1129, L1108, L1151 ); 
   and2 U2351 ( L902, L929, L1002 ); 
   inv U2352 ( L929, L933 ); 
   and3 U2353 ( L1221, L1226, L1287, L1308 ); 
   and3 U2354 ( L1217, L1230, L1291, L1311 ); 
   and3 U2355 ( L1244, L1249, L1295, L1314 ); 
   and3 U2356 ( L1240, L1253, L1299, L1317 ); 
   and3 U2357 ( L1267, L1272, L1303, L1320 ); 
   and3 U2358 ( L1263, L1276, L1307, L1323 ); 
   inv U2359 ( L1726, L1730 ); 
   and2 U2360 ( L1702, L1726, L1789 ); 
   and2 U2361 ( L1957, L1935, L1981 ); 
   inv U2362 ( L5817, L5823 ); 
   nand2 U2363 ( L5817, L5824, L1986 ); 
   inv U2364 ( L5825, L5831 ); 
   nand2 U2365 ( L5825, L5832, L1989 ); 
   inv U2366 ( L5833, L5839 ); 
   nand2 U2367 ( L5833, L5840, L1993 ); 
   inv U2368 ( L5841, L5847 ); 
   nand2 U2369 ( L5841, L5848, L1996 ); 
   nand2 U2370 ( L5849, L5856, L2000 ); 
   nand2 U2371 ( L5857, L5864, L2004 ); 
   or4 U2372 ( L2351, L2492, L2493, L2494, L2495 ); 
   or5 U2373 ( L2417, L2511, L2512, L2513, L2514, L2515 ); 
   or4 U2374 ( L2597, L2754, L2755, L2756, L2757 ); 
   or2 U2375 ( L2629, L2767, L2768 ); 
   or5 U2376 ( L2652, L2776, L2777, L2778, L2779, L2780 ); 
   or2 U2377 ( L2715, L2800, L2801 ); 
   or2 U2378 ( L3028, L3045, L3046 ); 
   or4 U2379 ( L3059, L3128, L3129, L3130, L3131 ); 
   or5 U2380 ( L3090, L3139, L3140, L3141, L3142, L3143 ); 
   inv U2381 ( L3235, L3238 ); 
   and2 U2382 ( L3216, L3235, L3258 ); 
   or4 U2383 ( L3292, L3434, L3435, L3436, L3437 ); 
   or5 U2384 ( L3362, L3449, L3450, L3451, L3452, L3453 ); 
   and3 U2385 ( L3508, L3513, L3574, L3595 ); 
   and3 U2386 ( L3504, L3517, L3578, L3598 ); 
   or4 U2387 ( L3853, L4007, L4008, L4009, L4010 ); 
   or2 U2388 ( L3885, L4016, L4017 ); 
   or5 U2389 ( L3908, L4024, L4025, L4026, L4027, L4028 ); 
   or2 U2390 ( L3971, L4047, L4048 ); 
   and3 U2391 ( L4230, L4235, L4266, L4283 ); 
   and3 U2392 ( L4226, L4239, L4270, L4286 ); 
   or4 U2393 ( L4297, L4361, L4362, L4363, L4364 ); 
   or5 U2394 ( L4324, L4372, L4373, L4374, L4375, L4376 ); 
   and3 U2395 ( L4535, L4540, L4601, L4622 ); 
   and3 U2396 ( L4531, L4544, L4605, L4625 ); 
   nand2 U2397 ( L4942, L4945, L4947 ); 
   nand2 U2398 ( L4983, L4986, L4988 ); 
   inv U2399 ( L5014, L5018 ); 
   nand2 U2400 ( L5014, L5017, L5019 ); 
   or2 U2401 ( L950, L956, L5024 ); 
   inv U2402 ( L5034, L5038 ); 
   inv U2403 ( L5102, L5106 ); 
   nand2 U2404 ( L5102, L5105, L5107 ); 
   inv U2405 ( L950, L5112 ); 
   inv U2406 ( L5122, L5126 ); 
   or2 U2407 ( L1715, L1749, L5468 ); 
   inv U2408 ( L5478, L5482 ); 
   inv U2409 ( L1715, L5526 ); 
   inv U2410 ( L5536, L5540 ); 
   inv U2411 ( L5584, L5588 ); 
   nand2 U2412 ( L5584, L5587, L5589 ); 
   or2 U2413 ( L1746, L1750, L5594 ); 
   inv U2414 ( L5604, L5608 ); 
   inv U2415 ( L5672, L5676 ); 
   nand2 U2416 ( L5672, L5675, L5677 ); 
   inv U2417 ( L1746, L5682 ); 
   inv U2418 ( L5692, L5696 ); 
   or4 U2419 ( L2366, L2500, L2501, L2502, L5937 ); 
   nor3 U2420 ( L2366, L2503, L2504, L5945 ); 
   or3 U2421 ( L2384, L2505, L2506, L5953 ); 
   nor2 U2422 ( L2384, L2507, L5961 ); 
   or4 U2423 ( L2612, L2762, L2763, L2764, L6070 ); 
   nor3 U2424 ( L2612, L2765, L2766, L6128 ); 
   nor3 U2425 ( L2693, L2798, L2799, L6264 ); 
   nor4 U2426 ( L2670, L2792, L2793, L2794, L6284 ); 
   nand2 U2427 ( L7348, L7351, L6360 ); 
   nand2 U2428 ( L7345, L7352, L6361 ); 
   or4 U2429 ( L3308, L3438, L3439, L3440, L6639 ); 
   nor3 U2430 ( L3308, L3441, L3442, L6647 ); 
   or3 U2431 ( L3327, L3443, L3444, L6655 ); 
   nor2 U2432 ( L3327, L3445, L6663 ); 
   nand2 U2433 ( L6812, L6815, L6817 ); 
   nand2 U2434 ( L6809, L6816, L6818 ); 
   nand2 U2435 ( L6822, L6825, L6827 ); 
   nand2 U2436 ( L6819, L6826, L6828 ); 
   or4 U2437 ( L3868, L4011, L4012, L4013, L6938 ); 
   nor3 U2438 ( L3868, L4014, L4015, L6996 ); 
   or4 U2439 ( L3949, L4042, L4043, L4044, L7044 ); 
   or5 U2440 ( L3926, L4035, L4036, L4037, L4038, L7064 ); 
   nor3 U2441 ( L3949, L4045, L4046, L7132 ); 
   nor4 U2442 ( L3926, L4039, L4040, L4041, L7152 ); 
   nand2 U2443 ( L7614, L7617, L7446 ); 
   nand2 U2444 ( L7611, L7618, L7447 ); 
   nand2 U2445 ( L7606, L7609, L7456 ); 
   nand2 U2446 ( L7603, L7610, L7457 ); 
   or2 U2447 ( L1117, L1151, L241 ); 
   or2 U2448 ( L908, L1002, L265 ); 
   nand2 U2449 ( L2003, L2004, L2005 ); 
   inv U2450 ( L4796, L4800 ); 
   inv U2451 ( L4804, L4808 ); 
   inv U2452 ( L4812, L4816 ); 
   inv U2453 ( L4820, L4824 ); 
   inv U2454 ( L4828, L4832 ); 
   inv U2455 ( L4844, L4848 ); 
   inv U2456 ( L4852, L4856 ); 
   inv U2457 ( L4860, L4864 ); 
   inv U2458 ( L4868, L4872 ); 
   nor2 U2459 ( L1308, L1309, L1310 ); 
   nor2 U2460 ( L1311, L1312, L1313 ); 
   nor2 U2461 ( L1314, L1315, L1316 ); 
   nor2 U2462 ( L1317, L1318, L1319 ); 
   nor2 U2463 ( L1320, L1321, L1322 ); 
   nor2 U2464 ( L1323, L1324, L1325 ); 
   inv U2465 ( L5388, L5392 ); 
   or2 U2466 ( L1708, L1789, L1790 ); 
   or2 U2467 ( L1941, L1981, L1982 ); 
   nand2 U2468 ( L5820, L5823, L1985 ); 
   nand2 U2469 ( L5828, L5831, L1988 ); 
   nand2 U2470 ( L5836, L5839, L1992 ); 
   nand2 U2471 ( L5844, L5847, L1995 ); 
   nand2 U2472 ( L1999, L2000, L2001 ); 
   inv U2473 ( L2487, L2491 ); 
   and5 U2474 ( L2420, L2472, L2436, L2409, L2454, L2508 ); 
   and5 U2475 ( L4526, L2472, L2436, L2454, L2420, L2522 ); 
   and4 U2476 ( L4526, L2472, L2436, L2454, L2526 ); 
   and3 U2477 ( L4526, L2472, L2454, L2529 ); 
   and2 U2478 ( L4526, L2472, L2531 ); 
   inv U2479 ( L5940, L5944 ); 
   inv U2480 ( L5948, L5952 ); 
   inv U2481 ( L5956, L5960 ); 
   inv U2482 ( L5964, L5968 ); 
   nand2 U2483 ( L5972, L5975, L2555 ); 
   inv U2484 ( L5972, L5976 ); 
   nand2 U2485 ( L5980, L5983, L2559 ); 
   inv U2486 ( L5980, L5984 ); 
   inv U2487 ( L2749, L2753 ); 
   and5 U2488 ( L2742, L2701, L2676, L2655, L2643, L2771 ); 
   and4 U2489 ( L2742, L2676, L2655, L2701, L2791 ); 
   and3 U2490 ( L2742, L2676, L2701, L2797 ); 
   and2 U2491 ( L2742, L2701, L2807 ); 
   inv U2492 ( L6110, L6114 ); 
   inv U2493 ( L6168, L6172 ); 
   inv U2494 ( L6246, L6250 ); 
   inv U2495 ( L6256, L6260 ); 
   inv U2496 ( L6342, L6346 ); 
   inv U2497 ( L6352, L6356 ); 
   inv U2498 ( L3123, L3127 ); 
   and2 U2499 ( L3123, L3136, L3156 ); 
   or2 U2500 ( L3223, L3258, L3259 ); 
   and2 U2501 ( L3431, L3446, L3466 ); 
   inv U2502 ( L6642, L6646 ); 
   inv U2503 ( L6650, L6654 ); 
   inv U2504 ( L6658, L6662 ); 
   inv U2505 ( L6666, L6670 ); 
   nand2 U2506 ( L6674, L6677, L3483 ); 
   inv U2507 ( L6674, L6678 ); 
   nand2 U2508 ( L6682, L6685, L3487 ); 
   inv U2509 ( L6682, L6686 ); 
   inv U2510 ( L3579, L3582 ); 
   inv U2511 ( L3583, L3586 ); 
   inv U2512 ( L3587, L3590 ); 
   inv U2513 ( L3591, L3594 ); 
   nor2 U2514 ( L3595, L3596, L3597 ); 
   nor2 U2515 ( L3598, L3599, L3600 ); 
   and3 U2516 ( L3536, L3527, L3579, L3602 ); 
   and3 U2517 ( L3540, L3531, L3583, L3605 ); 
   and3 U2518 ( L3559, L3550, L3587, L3608 ); 
   and3 U2519 ( L3563, L3554, L3591, L3611 ); 
   inv U2520 ( L4020, L4023 ); 
   inv U2521 ( L6978, L6982 ); 
   inv U2522 ( L7036, L7040 ); 
   inv U2523 ( L7114, L7118 ); 
   inv U2524 ( L7124, L7128 ); 
   and2 U2525 ( L4004, L4020, L4089 ); 
   inv U2526 ( L4247, L4250 ); 
   inv U2527 ( L4251, L4254 ); 
   inv U2528 ( L4255, L4258 ); 
   inv U2529 ( L4259, L4262 ); 
   and3 U2530 ( L4189, L4180, L4247, L4272 ); 
   and3 U2531 ( L4193, L4184, L4251, L4275 ); 
   and3 U2532 ( L4212, L4203, L4255, L4278 ); 
   and3 U2533 ( L4216, L4207, L4259, L4281 ); 
   nor2 U2534 ( L4283, L4284, L4285 ); 
   nor2 U2535 ( L4286, L4287, L4288 ); 
   inv U2536 ( L4356, L4360 ); 
   nand2 U2537 ( L4369, L89, L4380 ); 
   and2 U2538 ( L4356, L4369, L4386 ); 
   inv U2539 ( L7438, L7442 ); 
   inv U2540 ( L4606, L4609 ); 
   inv U2541 ( L4610, L4613 ); 
   inv U2542 ( L4614, L4617 ); 
   inv U2543 ( L4618, L4621 ); 
   nor2 U2544 ( L4622, L4623, L4624 ); 
   nor2 U2545 ( L4625, L4626, L4627 ); 
   and3 U2546 ( L4563, L4554, L4606, L4629 ); 
   and3 U2547 ( L4567, L4558, L4610, L4632 ); 
   and3 U2548 ( L4586, L4577, L4614, L4635 ); 
   and3 U2549 ( L4590, L4581, L4618, L4638 ); 
   buffer U2550 ( L2472, L4836 ); 
   nand2 U2551 ( L4947, L4948, L4949 ); 
   nand2 U2552 ( L4988, L4989, L4990 ); 
   nand2 U2553 ( L5011, L5018, L5020 ); 
   nand2 U2554 ( L5099, L5106, L5108 ); 
   nand2 U2555 ( L5581, L5588, L5590 ); 
   nand2 U2556 ( L5669, L5676, L5678 ); 
   inv U2557 ( L6080, L6084 ); 
   inv U2558 ( L6090, L6094 ); 
   inv U2559 ( L6100, L6104 ); 
   inv U2560 ( L6138, L6142 ); 
   inv U2561 ( L6148, L6152 ); 
   inv U2562 ( L6158, L6162 ); 
   buffer U2563 ( L2742, L6206 ); 
   inv U2564 ( L6216, L6220 ); 
   inv U2565 ( L6226, L6230 ); 
   inv U2566 ( L6236, L6240 ); 
   inv U2567 ( L6324, L6328 ); 
   buffer U2568 ( L2742, L6294 ); 
   inv U2569 ( L6304, L6308 ); 
   inv U2570 ( L6314, L6318 ); 
   nand2 U2571 ( L6360, L6361, L6362 ); 
   nand2 U2572 ( L6817, L6818, L6840 ); 
   nand2 U2573 ( L6827, L6828, L6848 ); 
   inv U2574 ( L6948, L6952 ); 
   inv U2575 ( L6958, L6962 ); 
   inv U2576 ( L6968, L6972 ); 
   inv U2577 ( L7006, L7010 ); 
   inv U2578 ( L7016, L7020 ); 
   inv U2579 ( L7026, L7030 ); 
   inv U2580 ( L7074, L7078 ); 
   inv U2581 ( L7084, L7088 ); 
   inv U2582 ( L7094, L7098 ); 
   inv U2583 ( L7104, L7108 ); 
   inv U2584 ( L7192, L7196 ); 
   inv U2585 ( L7162, L7166 ); 
   inv U2586 ( L7172, L7176 ); 
   inv U2587 ( L7182, L7186 ); 
   nand2 U2588 ( L7446, L7447, L7448 ); 
   nand2 U2589 ( L7456, L7457, L7458 ); 
   and2 U2590 ( L3046, L3249, L254 ); 
   and2 U2591 ( L3046, L3249, L260 ); 
   nand2 U2592 ( L1985, L1986, L1987 ); 
   nand2 U2593 ( L1992, L1993, L1994 ); 
   inv U2594 ( L2001, L2002 ); 
   and2 U2595 ( L933, L924, L962 ); 
   and2 U2596 ( L1730, L1721, L1751 ); 
   nand2 U2597 ( L1988, L1989, L1990 ); 
   nand2 U2598 ( L1995, L1996, L1997 ); 
   inv U2599 ( L2495, L2499 ); 
   and2 U2600 ( L2515, L2487, L2536 ); 
   inv U2601 ( L5937, L5943 ); 
   nand2 U2602 ( L5937, L5944, L2542 ); 
   inv U2603 ( L5945, L5951 ); 
   nand2 U2604 ( L5945, L5952, L2545 ); 
   inv U2605 ( L5953, L5959 ); 
   nand2 U2606 ( L5953, L5960, L2549 ); 
   inv U2607 ( L5961, L5967 ); 
   nand2 U2608 ( L5961, L5968, L2552 ); 
   nand2 U2609 ( L5969, L5976, L2556 ); 
   nand2 U2610 ( L5977, L5984, L2560 ); 
   inv U2611 ( L2757, L2761 ); 
   inv U2612 ( L2780, L2784 ); 
   and2 U2613 ( L2749, L2780, L2853 ); 
   inv U2614 ( L3131, L3135 ); 
   inv U2615 ( L3143, L3146 ); 
   and2 U2616 ( L3123, L3143, L3163 ); 
   and2 U2617 ( L3453, L3431, L3467 ); 
   inv U2618 ( L6639, L6645 ); 
   nand2 U2619 ( L6639, L6646, L3470 ); 
   inv U2620 ( L6647, L6653 ); 
   nand2 U2621 ( L6647, L6654, L3473 ); 
   inv U2622 ( L6655, L6661 ); 
   nand2 U2623 ( L6655, L6662, L3477 ); 
   inv U2624 ( L6663, L6669 ); 
   nand2 U2625 ( L6663, L6670, L3480 ); 
   nand2 U2626 ( L6671, L6678, L3484 ); 
   nand2 U2627 ( L6679, L6686, L3488 ); 
   and3 U2628 ( L3531, L3536, L3582, L3601 ); 
   and3 U2629 ( L3527, L3540, L3586, L3604 ); 
   and3 U2630 ( L3554, L3559, L3590, L3607 ); 
   and3 U2631 ( L3550, L3563, L3594, L3610 ); 
   inv U2632 ( L4028, L4032 ); 
   and2 U2633 ( L4004, L4028, L4090 ); 
   and3 U2634 ( L4184, L4189, L4250, L4271 ); 
   and3 U2635 ( L4180, L4193, L4254, L4274 ); 
   and3 U2636 ( L4207, L4212, L4258, L4277 ); 
   and3 U2637 ( L4203, L4216, L4262, L4280 ); 
   inv U2638 ( L4364, L4368 ); 
   inv U2639 ( L4376, L4379 ); 
   and2 U2640 ( L4356, L4376, L4387 ); 
   and3 U2641 ( L4558, L4563, L4609, L4628 ); 
   and3 U2642 ( L4554, L4567, L4613, L4631 ); 
   and3 U2643 ( L4581, L4586, L4617, L4634 ); 
   and3 U2644 ( L4577, L4590, L4621, L4637 ); 
   or5 U2645 ( L2431, L2518, L2519, L2520, L2522, L4841 ); 
   or4 U2646 ( L2448, L2523, L2524, L2526, L4849 ); 
   or3 U2647 ( L2465, L2527, L2529, L4857 ); 
   or2 U2648 ( L2481, L2531, L4865 ); 
   nand2 U2649 ( L5019, L5020, L5021 ); 
   inv U2650 ( L5024, L5028 ); 
   nand2 U2651 ( L5107, L5108, L5109 ); 
   inv U2652 ( L5112, L5116 ); 
   nand2 U2653 ( L1313, L1310, L5369 ); 
   nand2 U2654 ( L1319, L1316, L5377 ); 
   nand2 U2655 ( L1325, L1322, L5385 ); 
   inv U2656 ( L5468, L5472 ); 
   nand2 U2657 ( L5468, L5471, L5473 ); 
   inv U2658 ( L5526, L5530 ); 
   nand2 U2659 ( L5526, L5529, L5531 ); 
   nand2 U2660 ( L5589, L5590, L5591 ); 
   inv U2661 ( L5594, L5598 ); 
   nand2 U2662 ( L5677, L5678, L5679 ); 
   inv U2663 ( L5682, L5686 ); 
   or2 U2664 ( L2768, L2804, L6060 ); 
   inv U2665 ( L6070, L6074 ); 
   inv U2666 ( L2768, L6118 ); 
   inv U2667 ( L6128, L6132 ); 
   or4 U2668 ( L2693, L2795, L2796, L2797, L6176 ); 
   or2 U2669 ( L2801, L2807, L6186 ); 
   or5 U2670 ( L2670, L2788, L2789, L2790, L2791, L6196 ); 
   inv U2671 ( L6264, L6268 ); 
   nand2 U2672 ( L6264, L6267, L6269 ); 
   inv U2673 ( L2801, L6274 ); 
   inv U2674 ( L6284, L6288 ); 
   nand2 U2675 ( L4288, L4285, L6337 ); 
   nand2 U2676 ( L3600, L3597, L6829 ); 
   or2 U2677 ( L4017, L4051, L6928 ); 
   inv U2678 ( L6938, L6942 ); 
   inv U2679 ( L4017, L6986 ); 
   inv U2680 ( L6996, L7000 ); 
   inv U2681 ( L7044, L7048 ); 
   nand2 U2682 ( L7044, L7047, L7049 ); 
   or2 U2683 ( L4048, L4052, L7054 ); 
   inv U2684 ( L7064, L7068 ); 
   inv U2685 ( L7132, L7136 ); 
   nand2 U2686 ( L7132, L7135, L7137 ); 
   inv U2687 ( L4048, L7142 ); 
   inv U2688 ( L7152, L7156 ); 
   nand2 U2689 ( L4627, L4624, L7433 ); 
   and2 U2690 ( L1982, L1146, L242 ); 
   nand2 U2691 ( L3135, L3127, L3151 ); 
   and5 U2692 ( L89, L4386, L3156, L3035, L3249, L257 ); 
   and5 U2693 ( L89, L4386, L3156, L3035, L3249, L263 ); 
   and2 U2694 ( L1790, L997, L266 ); 
   inv U2695 ( L1990, L1991 ); 
   inv U2696 ( L1997, L1998 ); 
   nand2 U2697 ( L3487, L3488, L3489 ); 
   nand2 U2698 ( L4836, L4839, L371 ); 
   inv U2699 ( L4836, L4840 ); 
   nand2 U2700 ( L2559, L2560, L2561 ); 
   and2 U2701 ( L2487, L2508, L2532 ); 
   or2 U2702 ( L2495, L2536, L2537 ); 
   nand2 U2703 ( L5940, L5943, L2541 ); 
   nand2 U2704 ( L5948, L5951, L2544 ); 
   nand2 U2705 ( L5956, L5959, L2548 ); 
   nand2 U2706 ( L5964, L5967, L2551 ); 
   nand2 U2707 ( L2555, L2556, L2557 ); 
   and2 U2708 ( L2508, L4526, L2563 ); 
   nand2 U2709 ( L2499, L2491, L2577 ); 
   inv U2710 ( L2771, L2775 ); 
   nand2 U2711 ( L2771, L4526, L2806 ); 
   nand2 U2712 ( L2761, L2753, L2808 ); 
   and2 U2713 ( L2749, L2771, L2852 ); 
   or2 U2714 ( L2757, L2853, L2854 ); 
   inv U2715 ( L6362, L6366 ); 
   nand2 U2716 ( L4368, L4360, L4381 ); 
   or2 U2717 ( L3131, L3163, L3164 ); 
   and4 U2718 ( L89, L4386, L3156, L3035, L3241 ); 
   or2 U2719 ( L3437, L3467, L3468 ); 
   nand2 U2720 ( L6642, L6645, L3469 ); 
   nand2 U2721 ( L6650, L6653, L3472 ); 
   nand2 U2722 ( L6658, L6661, L3476 ); 
   nand2 U2723 ( L6666, L6669, L3479 ); 
   nand2 U2724 ( L3483, L3484, L3485 ); 
   nor2 U2725 ( L3601, L3602, L3603 ); 
   nor2 U2726 ( L3604, L3605, L3606 ); 
   nor2 U2727 ( L3607, L3608, L3609 ); 
   nor2 U2728 ( L3610, L3611, L3612 ); 
   inv U2729 ( L6840, L6844 ); 
   inv U2730 ( L6848, L6852 ); 
   or2 U2731 ( L4010, L4090, L4091 ); 
   nor2 U2732 ( L4271, L4272, L4273 ); 
   nor2 U2733 ( L4274, L4275, L4276 ); 
   nor2 U2734 ( L4277, L4278, L4279 ); 
   nor2 U2735 ( L4280, L4281, L4282 ); 
   and2 U2736 ( L4379, L4380, L4382 ); 
   or2 U2737 ( L4364, L4387, L4388 ); 
   inv U2738 ( L7448, L7452 ); 
   inv U2739 ( L7458, L7462 ); 
   nor2 U2740 ( L4628, L4629, L4630 ); 
   nor2 U2741 ( L4631, L4632, L4633 ); 
   nor2 U2742 ( L4634, L4635, L4636 ); 
   nor2 U2743 ( L4637, L4638, L4639 ); 
   inv U2744 ( L4949, L4955 ); 
   nand2 U2745 ( L4949, L4956, L4958 ); 
   inv U2746 ( L4990, L4996 ); 
   nand2 U2747 ( L4990, L4997, L4999 ); 
   nand2 U2748 ( L5465, L5472, L5474 ); 
   nand2 U2749 ( L5523, L5530, L5532 ); 
   inv U2750 ( L6206, L6210 ); 
   nand2 U2751 ( L6261, L6268, L6270 ); 
   inv U2752 ( L6294, L6298 ); 
   nand2 U2753 ( L7041, L7048, L7050 ); 
   nand2 U2754 ( L7129, L7136, L7138 ); 
   nand2 U2755 ( L3469, L3470, L3471 ); 
   nand2 U2756 ( L3476, L3477, L3478 ); 
   inv U2757 ( L3485, L3486 ); 
   nand2 U2758 ( L4833, L4840, L372 ); 
   nand2 U2759 ( L2541, L2542, L2543 ); 
   nand2 U2760 ( L2548, L2549, L2550 ); 
   inv U2761 ( L2557, L2558 ); 
   inv U2762 ( L4841, L4847 ); 
   nand2 U2763 ( L4841, L4848, L387 ); 
   inv U2764 ( L4849, L4855 ); 
   nand2 U2765 ( L4849, L4856, L390 ); 
   inv U2766 ( L4857, L4863 ); 
   nand2 U2767 ( L4857, L4864, L393 ); 
   inv U2768 ( L4865, L4871 ); 
   nand2 U2769 ( L4865, L4872, L396 ); 
   inv U2770 ( L962, L965 ); 
   inv U2771 ( L5369, L5375 ); 
   nand2 U2772 ( L5369, L5376, L1327 ); 
   inv U2773 ( L5377, L5383 ); 
   nand2 U2774 ( L5377, L5384, L1330 ); 
   inv U2775 ( L5385, L5391 ); 
   nand2 U2776 ( L5385, L5392, L1333 ); 
   inv U2777 ( L1751, L1754 ); 
   nand2 U2778 ( L2544, L2545, L2546 ); 
   nand2 U2779 ( L2551, L2552, L2553 ); 
   or2 U2780 ( L2515, L2563, L2564 ); 
   and2 U2781 ( L2784, L2806, L2809 ); 
   and2 U2782 ( L2784, L2775, L2813 ); 
   inv U2783 ( L6337, L6345 ); 
   nand2 U2784 ( L6337, L6346, L2860 ); 
   nand2 U2785 ( L3472, L3473, L3474 ); 
   nand2 U2786 ( L3479, L3480, L3481 ); 
   inv U2787 ( L6829, L6835 ); 
   nand2 U2788 ( L6829, L6836, L3614 ); 
   and2 U2789 ( L4032, L4023, L4053 ); 
   inv U2790 ( L7433, L7441 ); 
   nand2 U2791 ( L7433, L7442, L4516 ); 
   nand2 U2792 ( L4952, L4955, L4957 ); 
   nand2 U2793 ( L4993, L4996, L4998 ); 
   inv U2794 ( L5021, L5027 ); 
   nand2 U2795 ( L5021, L5028, L5030 ); 
   inv U2796 ( L5109, L5115 ); 
   nand2 U2797 ( L5109, L5116, L5118 ); 
   nand2 U2798 ( L5473, L5474, L5475 ); 
   nand2 U2799 ( L5531, L5532, L5533 ); 
   inv U2800 ( L5591, L5597 ); 
   nand2 U2801 ( L5591, L5598, L5600 ); 
   inv U2802 ( L5679, L5685 ); 
   nand2 U2803 ( L5679, L5686, L5688 ); 
   inv U2804 ( L6060, L6064 ); 
   nand2 U2805 ( L6060, L6063, L6065 ); 
   inv U2806 ( L6118, L6122 ); 
   nand2 U2807 ( L6118, L6121, L6123 ); 
   inv U2808 ( L6176, L6180 ); 
   nand2 U2809 ( L6176, L6179, L6181 ); 
   inv U2810 ( L6186, L6190 ); 
   inv U2811 ( L6196, L6200 ); 
   nand2 U2812 ( L6269, L6270, L6271 ); 
   inv U2813 ( L6274, L6278 ); 
   nand2 U2814 ( L4276, L4273, L6347 ); 
   nand2 U2815 ( L4282, L4279, L6357 ); 
   nand2 U2816 ( L3606, L3603, L6837 ); 
   nand2 U2817 ( L3612, L3609, L6845 ); 
   inv U2818 ( L6928, L6932 ); 
   nand2 U2819 ( L6928, L6931, L6933 ); 
   inv U2820 ( L6986, L6990 ); 
   nand2 U2821 ( L6986, L6989, L6991 ); 
   nand2 U2822 ( L7049, L7050, L7051 ); 
   inv U2823 ( L7054, L7058 ); 
   nand2 U2824 ( L7137, L7138, L7139 ); 
   inv U2825 ( L7142, L7146 ); 
   nand2 U2826 ( L4639, L4636, L7443 ); 
   nand2 U2827 ( L4633, L4630, L7453 ); 
   and3 U2828 ( L3468, L1974, L1146, L243 ); 
   and4 U2829 ( L2537, L3466, L1974, L1146, L244 ); 
   and5 U2830 ( L4526, L2532, L3466, L1974, L1146, L245 ); 
   and3 U2831 ( L3164, L3035, L3249, L255 ); 
   and4 U2832 ( L4388, L3156, L3035, L3249, L256 ); 
   and3 U2833 ( L3164, L3035, L3249, L261 ); 
   and4 U2834 ( L4388, L3156, L3035, L3249, L262 ); 
   and3 U2835 ( L4091, L1788, L997, L267 ); 
   and4 U2836 ( L2854, L4089, L1788, L997, L268 ); 
   and5 U2837 ( L4526, L2852, L4089, L1788, L997, L269 ); 
   inv U2838 ( L3474, L3475 ); 
   inv U2839 ( L3481, L3482 ); 
   nand2 U2840 ( L371, L372, L373 ); 
   inv U2841 ( L2546, L2547 ); 
   inv U2842 ( L2553, L2554 ); 
   nand2 U2843 ( L4844, L4847, L386 ); 
   nand2 U2844 ( L4852, L4855, L389 ); 
   nand2 U2845 ( L4860, L4863, L392 ); 
   nand2 U2846 ( L4868, L4871, L395 ); 
   nand2 U2847 ( L5372, L5375, L1326 ); 
   nand2 U2848 ( L5380, L5383, L1329 ); 
   nand2 U2849 ( L5388, L5391, L1332 ); 
   and2 U2850 ( L4091, L1788, L1436 ); 
   and3 U2851 ( L2854, L4089, L1788, L1440 ); 
   and4 U2852 ( L4526, L2852, L4089, L1788, L1445 ); 
   and2 U2853 ( L2854, L4089, L1450 ); 
   and3 U2854 ( L4526, L2852, L4089, L1454 ); 
   nand2 U2855 ( L6342, L6345, L2859 ); 
   inv U2856 ( L4382, L4385 ); 
   and2 U2857 ( L4382, L4364, L3148 ); 
   and2 U2858 ( L3164, L3035, L3239 ); 
   and3 U2859 ( L4388, L3156, L3035, L3240 ); 
   and2 U2860 ( L3468, L1974, L3265 ); 
   and3 U2861 ( L2537, L3466, L1974, L3267 ); 
   and4 U2862 ( L4526, L2532, L3466, L1974, L3270 ); 
   and2 U2863 ( L2537, L3466, L3274 ); 
   and3 U2864 ( L4526, L2532, L3466, L3277 ); 
   nand2 U2865 ( L6832, L6835, L3613 ); 
   nand2 U2866 ( L7438, L7441, L4515 ); 
   nand2 U2867 ( L4957, L4958, L4959 ); 
   nand2 U2868 ( L4998, L4999, L5000 ); 
   nand2 U2869 ( L5024, L5027, L5029 ); 
   nand2 U2870 ( L5112, L5115, L5117 ); 
   nand2 U2871 ( L5594, L5597, L5599 ); 
   nand2 U2872 ( L5682, L5685, L5687 ); 
   nand2 U2873 ( L6057, L6064, L6066 ); 
   nand2 U2874 ( L6115, L6122, L6124 ); 
   nand2 U2875 ( L6173, L6180, L6182 ); 
   nand2 U2876 ( L6925, L6932, L6934 ); 
   nand2 U2877 ( L6983, L6990, L6992 ); 
   or5 U2878 ( L241, L242, L243, L244, L245, L246 ); 
   or5 U2879 ( L3259, L254, L255, L256, L257, L258 ); 
   or5 U2880 ( L3259, L260, L261, L262, L263, L264 ); 
   or5 U2881 ( L265, L266, L267, L268, L269, L270 ); 
   and2 U2882 ( L2564, L2543, L375 ); 
   and2 U2883 ( L2564, L2550, L378 ); 
   and2 U2884 ( L2564, L2558, L381 ); 
   and2 U2885 ( L2564, L2406, L384 ); 
   nand2 U2886 ( L386, L387, L388 ); 
   nand2 U2887 ( L389, L390, L391 ); 
   nand2 U2888 ( L392, L393, L394 ); 
   nand2 U2889 ( L395, L396, L397 ); 
   nand2 U2890 ( L1326, L1327, L1328 ); 
   nand2 U2891 ( L1329, L1330, L1331 ); 
   nand2 U2892 ( L1332, L1333, L1334 ); 
   or4 U2893 ( L1790, L1436, L1440, L1445, L1447 ); 
   or3 U2894 ( L4091, L1450, L1454, L1766 ); 
   inv U2895 ( L2564, L2571 ); 
   and2 U2896 ( L2577, L2564, L2579 ); 
   inv U2897 ( L2809, L2812 ); 
   inv U2898 ( L2813, L2816 ); 
   and2 U2899 ( L2809, L2757, L2851 ); 
   nand2 U2900 ( L2859, L2860, L2861 ); 
   inv U2901 ( L6347, L6355 ); 
   nand2 U2902 ( L6347, L6356, L2863 ); 
   inv U2903 ( L6357, L6365 ); 
   nand2 U2904 ( L6357, L6366, L2866 ); 
   and2 U2905 ( L4381, L4385, L3147 ); 
   or4 U2906 ( L3046, L3239, L3240, L3241, L3242 ); 
   or4 U2907 ( L1982, L3265, L3267, L3270, L3271 ); 
   or3 U2908 ( L3468, L3274, L3277, L3279 ); 
   nand2 U2909 ( L3613, L3614, L3615 ); 
   inv U2910 ( L6837, L6843 ); 
   nand2 U2911 ( L6837, L6844, L3617 ); 
   inv U2912 ( L6845, L6851 ); 
   nand2 U2913 ( L6845, L6852, L3620 ); 
   inv U2914 ( L4053, L4056 ); 
   nand2 U2915 ( L4515, L4516, L4517 ); 
   inv U2916 ( L7443, L7451 ); 
   nand2 U2917 ( L7443, L7452, L4519 ); 
   inv U2918 ( L7453, L7461 ); 
   nand2 U2919 ( L7453, L7462, L4522 ); 
   nand2 U2920 ( L5029, L5030, L5031 ); 
   nand2 U2921 ( L5117, L5118, L5119 ); 
   inv U2922 ( L5475, L5481 ); 
   nand2 U2923 ( L5475, L5482, L5484 ); 
   inv U2924 ( L5533, L5539 ); 
   nand2 U2925 ( L5533, L5540, L5542 ); 
   nand2 U2926 ( L5599, L5600, L5601 ); 
   nand2 U2927 ( L5687, L5688, L5689 ); 
   nand2 U2928 ( L6065, L6066, L6067 ); 
   nand2 U2929 ( L6123, L6124, L6125 ); 
   nand2 U2930 ( L6181, L6182, L6183 ); 
   inv U2931 ( L6271, L6277 ); 
   nand2 U2932 ( L6271, L6278, L6280 ); 
   nand2 U2933 ( L6933, L6934, L6935 ); 
   nand2 U2934 ( L6991, L6992, L6993 ); 
   inv U2935 ( L7051, L7057 ); 
   nand2 U2936 ( L7051, L7058, L7060 ); 
   inv U2937 ( L7139, L7145 ); 
   nand2 U2938 ( L7139, L7146, L7148 ); 
   nand2 U2939 ( L4959, L4966, L4968 ); 
   nand2 U2940 ( L5000, L5007, L5009 ); 
   and2 U2941 ( L2808, L2812, L2850 ); 
   nand2 U2942 ( L6352, L6355, L2862 ); 
   nand2 U2943 ( L6362, L6365, L2865 ); 
   or2 U2944 ( L3147, L3148, L3149 ); 
   nand2 U2945 ( L3228, L3242, L3243 ); 
   nand2 U2946 ( L6840, L6843, L3616 ); 
   nand2 U2947 ( L6848, L6851, L3619 ); 
   nand2 U2948 ( L7448, L7451, L4518 ); 
   nand2 U2949 ( L7458, L7461, L4521 ); 
   inv U2950 ( L4959, L4965 ); 
   inv U2951 ( L5000, L5006 ); 
   nand2 U2952 ( L5478, L5481, L5483 ); 
   nand2 U2953 ( L5536, L5539, L5541 ); 
   nand2 U2954 ( L6274, L6277, L6279 ); 
   nand2 U2955 ( L7054, L7057, L7059 ); 
   nand2 U2956 ( L7142, L7145, L7147 ); 
   and2 U2957 ( L2547, L2571, L374 ); 
   and2 U2958 ( L2554, L2571, L377 ); 
   and2 U2959 ( L2561, L2571, L380 ); 
   and2 U2960 ( L2400, L2571, L383 ); 
   nand2 U2961 ( L920, L1447, L955 ); 
   nand2 U2962 ( L4962, L4965, L4967 ); 
   nand2 U2963 ( L5003, L5006, L5008 ); 
   buffer U2964 ( L1447, L975 ); 
   and5 U2965 ( L3271, L1093, L1055, L1074, L1038, L1136 ); 
   and4 U2966 ( L3271, L1093, L1055, L1074, L1140 ); 
   and3 U2967 ( L3271, L1093, L1074, L1143 ); 
   and2 U2968 ( L3271, L1093, L1145 ); 
   and2 U2969 ( L1122, L3271, L1160 ); 
   inv U2970 ( L1766, L1771 ); 
   and5 U2971 ( L3279, L1921, L1885, L1903, L1869, L1964 ); 
   and4 U2972 ( L3279, L1921, L1885, L1903, L1968 ); 
   and3 U2973 ( L3279, L1921, L1903, L1971 ); 
   and2 U2974 ( L3279, L1921, L1973 ); 
   and2 U2975 ( L1950, L3279, L2007 ); 
   and2 U2976 ( L2495, L2571, L2578 ); 
   nand2 U2977 ( L2862, L2863, L2864 ); 
   nand2 U2978 ( L2865, L2866, L2867 ); 
   nand2 U2979 ( L3136, L3149, L3150 ); 
   and2 U2980 ( L3238, L3243, L3245 ); 
   nand2 U2981 ( L3616, L3617, L3618 ); 
   nand2 U2982 ( L3619, L3620, L3621 ); 
   or2 U2983 ( L2850, L2851, L4067 ); 
   nand2 U2984 ( L4518, L4519, L4520 ); 
   nand2 U2985 ( L4521, L4522, L4523 ); 
   buffer U2986 ( L3279, L4713 ); 
   buffer U2987 ( L3271, L4753 ); 
   inv U2988 ( L5031, L5037 ); 
   nand2 U2989 ( L5031, L5038, L5040 ); 
   inv U2990 ( L5119, L5125 ); 
   nand2 U2991 ( L5119, L5126, L5128 ); 
   nand2 U2992 ( L5483, L5484, L5485 ); 
   nand2 U2993 ( L5541, L5542, L5543 ); 
   inv U2994 ( L5601, L5607 ); 
   nand2 U2995 ( L5601, L5608, L5610 ); 
   inv U2996 ( L5689, L5695 ); 
   nand2 U2997 ( L5689, L5696, L5698 ); 
   inv U2998 ( L6067, L6073 ); 
   nand2 U2999 ( L6067, L6074, L6076 ); 
   inv U3000 ( L6125, L6131 ); 
   nand2 U3001 ( L6125, L6132, L6134 ); 
   inv U3002 ( L6183, L6189 ); 
   nand2 U3003 ( L6183, L6190, L6192 ); 
   nand2 U3004 ( L6279, L6280, L6281 ); 
   inv U3005 ( L6935, L6941 ); 
   nand2 U3006 ( L6935, L6942, L6944 ); 
   inv U3007 ( L6993, L6999 ); 
   nand2 U3008 ( L6993, L7000, L7002 ); 
   nand2 U3009 ( L7059, L7060, L7061 ); 
   nand2 U3010 ( L7147, L7148, L7149 ); 
   or2 U3011 ( L374, L375, L376 ); 
   or2 U3012 ( L377, L378, L379 ); 
   or2 U3013 ( L380, L381, L382 ); 
   or2 U3014 ( L383, L384, L385 ); 
   and2 U3015 ( L933, L955, L958 ); 
   nand2 U3016 ( L4967, L4968, L967 ); 
   nand2 U3017 ( L5008, L5009, L971 ); 
   or2 U3018 ( L1129, L1160, L1161 ); 
   or2 U3019 ( L1957, L2007, L2008 ); 
   or2 U3020 ( L2578, L2579, L2580 ); 
   and4 U3021 ( L1331, L2861, L2864, L2867, L2868 ); 
   and2 U3022 ( L3146, L3150, L3152 ); 
   and4 U3023 ( L1328, L1334, L3618, L3621, L4443 ); 
   and4 U3024 ( L3615, L4517, L4520, L4523, L4524 ); 
   or5 U3025 ( L1880, L1960, L1961, L1962, L1964, L4721 ); 
   or4 U3026 ( L1897, L1965, L1966, L1968, L4729 ); 
   or3 U3027 ( L1914, L1969, L1971, L4737 ); 
   or2 U3028 ( L1929, L1973, L4745 ); 
   or5 U3029 ( L1050, L1132, L1133, L1134, L1136, L4761 ); 
   or4 U3030 ( L1068, L1137, L1138, L1140, L4769 ); 
   or3 U3031 ( L1086, L1141, L1143, L4777 ); 
   or2 U3032 ( L1102, L1145, L4785 ); 
   nand2 U3033 ( L5034, L5037, L5039 ); 
   nand2 U3034 ( L5122, L5125, L5127 ); 
   nand2 U3035 ( L5604, L5607, L5609 ); 
   nand2 U3036 ( L5692, L5695, L5697 ); 
   nand2 U3037 ( L6070, L6073, L6075 ); 
   nand2 U3038 ( L6128, L6131, L6133 ); 
   nand2 U3039 ( L6186, L6189, L6191 ); 
   nand2 U3040 ( L6938, L6941, L6943 ); 
   nand2 U3041 ( L6996, L6999, L7001 ); 
   inv U3042 ( L3245, L3248 ); 
   and2 U3043 ( L3245, L3223, L248 ); 
   inv U3044 ( L4713, L4719 ); 
   nand2 U3045 ( L4713, L4720, L294 ); 
   inv U3046 ( L4753, L4759 ); 
   nand2 U3047 ( L4753, L4760, L323 ); 
   inv U3048 ( L975, L980 ); 
   inv U3049 ( L4067, L4072 ); 
   nand2 U3050 ( L5039, L5040, L5041 ); 
   nand2 U3051 ( L5127, L5128, L5129 ); 
   inv U3052 ( L5485, L5491 ); 
   nand2 U3053 ( L5485, L5492, L5494 ); 
   inv U3054 ( L5543, L5549 ); 
   nand2 U3055 ( L5543, L5550, L5552 ); 
   nand2 U3056 ( L5609, L5610, L5611 ); 
   nand2 U3057 ( L5697, L5698, L5699 ); 
   nand2 U3058 ( L6075, L6076, L6077 ); 
   nand2 U3059 ( L6133, L6134, L6135 ); 
   nand2 U3060 ( L6191, L6192, L6193 ); 
   inv U3061 ( L6281, L6287 ); 
   nand2 U3062 ( L6281, L6288, L6290 ); 
   nand2 U3063 ( L6943, L6944, L6945 ); 
   nand2 U3064 ( L7001, L7002, L7003 ); 
   inv U3065 ( L7061, L7067 ); 
   nand2 U3066 ( L7061, L7068, L7070 ); 
   inv U3067 ( L7149, L7155 ); 
   nand2 U3068 ( L7149, L7156, L7158 ); 
   and2 U3069 ( L3244, L3248, L247 ); 
   inv U3070 ( L3152, L3155 ); 
   and2 U3071 ( L3152, L3131, L251 ); 
   and2 U3072 ( L1176, L1161, L272 ); 
   inv U3073 ( L958, L961 ); 
   and2 U3074 ( L958, L908, L275 ); 
   nand2 U3075 ( L4716, L4719, L293 ); 
   and2 U3076 ( L2008, L1987, L297 ); 
   and2 U3077 ( L2008, L1994, L300 ); 
   and2 U3078 ( L2008, L2002, L303 ); 
   and2 U3079 ( L2008, L1856, L306 ); 
   inv U3080 ( L4721, L4727 ); 
   nand2 U3081 ( L4721, L4728, L309 ); 
   inv U3082 ( L4729, L4735 ); 
   nand2 U3083 ( L4729, L4736, L312 ); 
   inv U3084 ( L4737, L4743 ); 
   nand2 U3085 ( L4737, L4744, L315 ); 
   inv U3086 ( L4745, L4751 ); 
   nand2 U3087 ( L4745, L4752, L318 ); 
   nand2 U3088 ( L4756, L4759, L322 ); 
   inv U3089 ( L4761, L4767 ); 
   nand2 U3090 ( L4761, L4768, L326 ); 
   inv U3091 ( L4769, L4775 ); 
   nand2 U3092 ( L4769, L4776, L329 ); 
   inv U3093 ( L4777, L4783 ); 
   nand2 U3094 ( L4777, L4784, L332 ); 
   inv U3095 ( L4785, L4791 ); 
   nand2 U3096 ( L4785, L4792, L335 ); 
   inv U3097 ( L4443, L412 ); 
   inv U3098 ( L4524, L414 ); 
   inv U3099 ( L2868, L416 ); 
   and3 U3100 ( L4443, L4524, L2868, L2881 ); 
   and3 U3101 ( L971, L962, L975, L993 ); 
   and3 U3102 ( L967, L965, L975, L994 ); 
   inv U3103 ( L1161, L1166 ); 
   and2 U3104 ( L1161, L1155, L1171 ); 
   and2 U3105 ( L1161, L1023, L1174 ); 
   inv U3106 ( L2008, L2014 ); 
   and5 U3107 ( L2580, L3417, L3381, L3399, L3365, L3459 ); 
   and4 U3108 ( L2580, L3417, L3381, L3399, L3462 ); 
   and3 U3109 ( L2580, L3417, L3399, L3464 ); 
   and2 U3110 ( L2580, L3417, L3465 ); 
   and2 U3111 ( L3446, L2580, L3490 ); 
   buffer U3112 ( L2580, L4793 ); 
   nand2 U3113 ( L5488, L5491, L5493 ); 
   nand2 U3114 ( L5546, L5549, L5551 ); 
   nand2 U3115 ( L6284, L6287, L6289 ); 
   nand2 U3116 ( L7064, L7067, L7069 ); 
   nand2 U3117 ( L7152, L7155, L7157 ); 
   or2 U3118 ( L247, L248, L249 ); 
   and2 U3119 ( L3151, L3155, L250 ); 
   and2 U3120 ( L957, L961, L274 ); 
   nand2 U3121 ( L293, L294, L295 ); 
   nand2 U3122 ( L4724, L4727, L308 ); 
   nand2 U3123 ( L4732, L4735, L311 ); 
   nand2 U3124 ( L4740, L4743, L314 ); 
   nand2 U3125 ( L4748, L4751, L317 ); 
   nand2 U3126 ( L322, L323, L324 ); 
   nand2 U3127 ( L4764, L4767, L325 ); 
   nand2 U3128 ( L4772, L4775, L328 ); 
   nand2 U3129 ( L4780, L4783, L331 ); 
   nand2 U3130 ( L4788, L4791, L334 ); 
   and3 U3131 ( L2876, L2878, L2881, L417 ); 
   and3 U3132 ( L971, L933, L980, L991 ); 
   and3 U3133 ( L967, L929, L980, L992 ); 
   or2 U3134 ( L3453, L3490, L3491 ); 
   or5 U3135 ( L3376, L3456, L3457, L3458, L3459, L4801 ); 
   or4 U3136 ( L3393, L3460, L3461, L3462, L4809 ); 
   or3 U3137 ( L3410, L3463, L3464, L4817 ); 
   or2 U3138 ( L3425, L3465, L4825 ); 
   inv U3139 ( L5041, L5047 ); 
   nand2 U3140 ( L5041, L5048, L5050 ); 
   inv U3141 ( L5129, L5135 ); 
   nand2 U3142 ( L5129, L5136, L5138 ); 
   nand2 U3143 ( L5493, L5494, L5495 ); 
   nand2 U3144 ( L5551, L5552, L5553 ); 
   inv U3145 ( L5611, L5617 ); 
   nand2 U3146 ( L5611, L5618, L5620 ); 
   inv U3147 ( L5699, L5705 ); 
   nand2 U3148 ( L5699, L5706, L5708 ); 
   inv U3149 ( L6077, L6083 ); 
   nand2 U3150 ( L6077, L6084, L6086 ); 
   inv U3151 ( L6135, L6141 ); 
   nand2 U3152 ( L6135, L6142, L6144 ); 
   inv U3153 ( L6193, L6199 ); 
   nand2 U3154 ( L6193, L6200, L6202 ); 
   nand2 U3155 ( L6289, L6290, L6291 ); 
   inv U3156 ( L6945, L6951 ); 
   nand2 U3157 ( L6945, L6952, L6954 ); 
   inv U3158 ( L7003, L7009 ); 
   nand2 U3159 ( L7003, L7010, L7012 ); 
   nand2 U3160 ( L7069, L7070, L7071 ); 
   nand2 U3161 ( L7157, L7158, L7159 ); 
   or2 U3162 ( L250, L251, L252 ); 
   and2 U3163 ( L1117, L1166, L271 ); 
   or2 U3164 ( L274, L275, L276 ); 
   and2 U3165 ( L1991, L2014, L296 ); 
   and2 U3166 ( L1998, L2014, L299 ); 
   and2 U3167 ( L2005, L2014, L302 ); 
   and2 U3168 ( L1850, L2014, L305 ); 
   nand2 U3169 ( L308, L309, L310 ); 
   nand2 U3170 ( L311, L312, L313 ); 
   nand2 U3171 ( L314, L315, L316 ); 
   nand2 U3172 ( L317, L318, L319 ); 
   nand2 U3173 ( L325, L326, L327 ); 
   nand2 U3174 ( L328, L329, L330 ); 
   nand2 U3175 ( L331, L332, L333 ); 
   nand2 U3176 ( L334, L335, L336 ); 
   inv U3177 ( L4793, L4799 ); 
   nand2 U3178 ( L4793, L4800, L343 ); 
   inv U3179 ( L417, L418 ); 
   and2 U3180 ( L1158, L1166, L1170 ); 
   and2 U3181 ( L1019, L1166, L1173 ); 
   nand2 U3182 ( L5044, L5047, L5049 ); 
   nand2 U3183 ( L5132, L5135, L5137 ); 
   or4 U3184 ( L991, L992, L993, L994, L5167 ); 
   nand2 U3185 ( L5614, L5617, L5619 ); 
   nand2 U3186 ( L5702, L5705, L5707 ); 
   nand2 U3187 ( L6080, L6083, L6085 ); 
   nand2 U3188 ( L6138, L6141, L6143 ); 
   nand2 U3189 ( L6196, L6199, L6201 ); 
   nand2 U3190 ( L6948, L6951, L6953 ); 
   nand2 U3191 ( L7006, L7009, L7011 ); 
   or2 U3192 ( L271, L272, L273 ); 
   or2 U3193 ( L296, L297, L298 ); 
   or2 U3194 ( L299, L300, L301 ); 
   or2 U3195 ( L302, L303, L304 ); 
   or2 U3196 ( L305, L306, L307 ); 
   nand2 U3197 ( L4796, L4799, L342 ); 
   and2 U3198 ( L3491, L3471, L346 ); 
   and2 U3199 ( L3491, L3478, L349 ); 
   and2 U3200 ( L3491, L3486, L352 ); 
   and2 U3201 ( L3491, L3350, L355 ); 
   inv U3202 ( L4801, L4807 ); 
   nand2 U3203 ( L4801, L4808, L358 ); 
   inv U3204 ( L4809, L4815 ); 
   nand2 U3205 ( L4809, L4816, L361 ); 
   inv U3206 ( L4817, L4823 ); 
   nand2 U3207 ( L4817, L4824, L364 ); 
   inv U3208 ( L4825, L4831 ); 
   nand2 U3209 ( L4825, L4832, L367 ); 
   or2 U3210 ( L1170, L1171, L1172 ); 
   or2 U3211 ( L1173, L1174, L1175 ); 
   inv U3212 ( L3491, L3497 ); 
   nand2 U3213 ( L5049, L5050, L5051 ); 
   nand2 U3214 ( L5137, L5138, L5139 ); 
   inv U3215 ( L5495, L5501 ); 
   nand2 U3216 ( L5495, L5502, L5504 ); 
   inv U3217 ( L5553, L5559 ); 
   nand2 U3218 ( L5553, L5560, L5562 ); 
   nand2 U3219 ( L5619, L5620, L5621 ); 
   nand2 U3220 ( L5707, L5708, L5709 ); 
   nand2 U3221 ( L6085, L6086, L6087 ); 
   nand2 U3222 ( L6143, L6144, L6145 ); 
   nand2 U3223 ( L6201, L6202, L6203 ); 
   inv U3224 ( L6291, L6297 ); 
   nand2 U3225 ( L6291, L6298, L6300 ); 
   nand2 U3226 ( L6953, L6954, L6955 ); 
   nand2 U3227 ( L7011, L7012, L7013 ); 
   inv U3228 ( L7071, L7077 ); 
   nand2 U3229 ( L7071, L7078, L7080 ); 
   inv U3230 ( L7159, L7165 ); 
   nand2 U3231 ( L7159, L7166, L7168 ); 
   nand2 U3232 ( L342, L343, L344 ); 
   nand2 U3233 ( L4804, L4807, L357 ); 
   nand2 U3234 ( L4812, L4815, L360 ); 
   nand2 U3235 ( L4820, L4823, L363 ); 
   nand2 U3236 ( L4828, L4831, L366 ); 
   inv U3237 ( L5167, L5173 ); 
   buffer U3238 ( L1172, L422 ); 
   buffer U3239 ( L1172, L469 ); 
   buffer U3240 ( L1175, L419 ); 
   buffer U3241 ( L1175, L471 ); 
   nand2 U3242 ( L5498, L5501, L5503 ); 
   nand2 U3243 ( L5556, L5559, L5561 ); 
   nand2 U3244 ( L6294, L6297, L6299 ); 
   nand2 U3245 ( L7074, L7077, L7079 ); 
   nand2 U3246 ( L7162, L7165, L7167 ); 
   and2 U3247 ( L3475, L3497, L345 ); 
   and2 U3248 ( L3482, L3497, L348 ); 
   and2 U3249 ( L3489, L3497, L351 ); 
   and2 U3250 ( L3344, L3497, L354 ); 
   nand2 U3251 ( L357, L358, L359 ); 
   nand2 U3252 ( L360, L361, L362 ); 
   nand2 U3253 ( L363, L364, L365 ); 
   nand2 U3254 ( L366, L367, L368 ); 
   inv U3255 ( L5051, L5057 ); 
   nand2 U3256 ( L5051, L5058, L5060 ); 
   inv U3257 ( L5139, L5145 ); 
   nand2 U3258 ( L5139, L5146, L5148 ); 
   nand2 U3259 ( L5503, L5504, L5505 ); 
   nand2 U3260 ( L5561, L5562, L5563 ); 
   inv U3261 ( L5621, L5627 ); 
   nand2 U3262 ( L5621, L5628, L5630 ); 
   inv U3263 ( L5709, L5715 ); 
   nand2 U3264 ( L5709, L5716, L5718 ); 
   inv U3265 ( L6087, L6093 ); 
   nand2 U3266 ( L6087, L6094, L6096 ); 
   inv U3267 ( L6145, L6151 ); 
   nand2 U3268 ( L6145, L6152, L6154 ); 
   inv U3269 ( L6203, L6209 ); 
   nand2 U3270 ( L6203, L6210, L6212 ); 
   nand2 U3271 ( L6299, L6300, L6301 ); 
   inv U3272 ( L6955, L6961 ); 
   nand2 U3273 ( L6955, L6962, L6964 ); 
   inv U3274 ( L7013, L7019 ); 
   nand2 U3275 ( L7013, L7020, L7022 ); 
   nand2 U3276 ( L7079, L7080, L7081 ); 
   nand2 U3277 ( L7167, L7168, L7169 ); 
   or2 U3278 ( L345, L346, L347 ); 
   or2 U3279 ( L348, L349, L350 ); 
   or2 U3280 ( L351, L352, L353 ); 
   or2 U3281 ( L354, L355, L356 ); 
   nand2 U3282 ( L5054, L5057, L5059 ); 
   nand2 U3283 ( L5142, L5145, L5147 ); 
   nand2 U3284 ( L5624, L5627, L5629 ); 
   nand2 U3285 ( L5712, L5715, L5717 ); 
   nand2 U3286 ( L6090, L6093, L6095 ); 
   nand2 U3287 ( L6148, L6151, L6153 ); 
   nand2 U3288 ( L6206, L6209, L6211 ); 
   nand2 U3289 ( L6958, L6961, L6963 ); 
   nand2 U3290 ( L7016, L7019, L7021 ); 
   nand2 U3291 ( L5059, L5060, L5061 ); 
   nand2 U3292 ( L5147, L5148, L5149 ); 
   inv U3293 ( L5505, L5511 ); 
   nand2 U3294 ( L5505, L5512, L5514 ); 
   inv U3295 ( L5563, L5569 ); 
   nand2 U3296 ( L5563, L5570, L5572 ); 
   nand2 U3297 ( L5629, L5630, L5631 ); 
   nand2 U3298 ( L5717, L5718, L5719 ); 
   nand2 U3299 ( L6095, L6096, L6097 ); 
   nand2 U3300 ( L6153, L6154, L6155 ); 
   nand2 U3301 ( L6211, L6212, L6213 ); 
   inv U3302 ( L6301, L6307 ); 
   nand2 U3303 ( L6301, L6308, L6310 ); 
   nand2 U3304 ( L6963, L6964, L6965 ); 
   nand2 U3305 ( L7021, L7022, L7023 ); 
   inv U3306 ( L7081, L7087 ); 
   nand2 U3307 ( L7081, L7088, L7090 ); 
   inv U3308 ( L7169, L7175 ); 
   nand2 U3309 ( L7169, L7176, L7178 ); 
   nand2 U3310 ( L5508, L5511, L5513 ); 
   nand2 U3311 ( L5566, L5569, L5571 ); 
   nand2 U3312 ( L6304, L6307, L6309 ); 
   nand2 U3313 ( L7084, L7087, L7089 ); 
   nand2 U3314 ( L7172, L7175, L7177 ); 
   inv U3315 ( L5061, L5067 ); 
   nand2 U3316 ( L5061, L5068, L5070 ); 
   inv U3317 ( L5149, L5155 ); 
   nand2 U3318 ( L5149, L5156, L5158 ); 
   nand2 U3319 ( L5513, L5514, L5515 ); 
   nand2 U3320 ( L5571, L5572, L5573 ); 
   inv U3321 ( L5631, L5637 ); 
   nand2 U3322 ( L5631, L5638, L5640 ); 
   inv U3323 ( L5719, L5725 ); 
   nand2 U3324 ( L5719, L5726, L5728 ); 
   inv U3325 ( L6097, L6103 ); 
   nand2 U3326 ( L6097, L6104, L6106 ); 
   inv U3327 ( L6155, L6161 ); 
   nand2 U3328 ( L6155, L6162, L6164 ); 
   inv U3329 ( L6213, L6219 ); 
   nand2 U3330 ( L6213, L6220, L6222 ); 
   nand2 U3331 ( L6309, L6310, L6311 ); 
   inv U3332 ( L6965, L6971 ); 
   nand2 U3333 ( L6965, L6972, L6974 ); 
   inv U3334 ( L7023, L7029 ); 
   nand2 U3335 ( L7023, L7030, L7032 ); 
   nand2 U3336 ( L7089, L7090, L7091 ); 
   nand2 U3337 ( L7177, L7178, L7179 ); 
   nand2 U3338 ( L5064, L5067, L5069 ); 
   nand2 U3339 ( L5152, L5155, L5157 ); 
   nand2 U3340 ( L5634, L5637, L5639 ); 
   nand2 U3341 ( L5722, L5725, L5727 ); 
   nand2 U3342 ( L6100, L6103, L6105 ); 
   nand2 U3343 ( L6158, L6161, L6163 ); 
   nand2 U3344 ( L6216, L6219, L6221 ); 
   nand2 U3345 ( L6968, L6971, L6973 ); 
   nand2 U3346 ( L7026, L7029, L7031 ); 
   inv U3347 ( L5515, L5521 ); 
   nand2 U3348 ( L5515, L5522, L1756 ); 
   inv U3349 ( L5573, L5579 ); 
   nand2 U3350 ( L5573, L5580, L1761 ); 
   nand2 U3351 ( L5069, L5070, L5071 ); 
   nand2 U3352 ( L5157, L5158, L5159 ); 
   nand2 U3353 ( L5639, L5640, L5641 ); 
   nand2 U3354 ( L5727, L5728, L5729 ); 
   nand2 U3355 ( L6105, L6106, L6107 ); 
   nand2 U3356 ( L6163, L6164, L6165 ); 
   nand2 U3357 ( L6221, L6222, L6223 ); 
   inv U3358 ( L6311, L6317 ); 
   nand2 U3359 ( L6311, L6318, L6320 ); 
   nand2 U3360 ( L6973, L6974, L6975 ); 
   nand2 U3361 ( L7031, L7032, L7033 ); 
   inv U3362 ( L7091, L7097 ); 
   nand2 U3363 ( L7091, L7098, L7100 ); 
   inv U3364 ( L7179, L7185 ); 
   nand2 U3365 ( L7179, L7186, L7188 ); 
   nand2 U3366 ( L5518, L5521, L1755 ); 
   nand2 U3367 ( L5576, L5579, L1760 ); 
   nand2 U3368 ( L6314, L6317, L6319 ); 
   nand2 U3369 ( L7094, L7097, L7099 ); 
   nand2 U3370 ( L7182, L7185, L7187 ); 
   nand2 U3371 ( L1755, L1756, L1757 ); 
   nand2 U3372 ( L1760, L1761, L1762 ); 
   inv U3373 ( L6107, L6113 ); 
   nand2 U3374 ( L6107, L6114, L2818 ); 
   inv U3375 ( L6165, L6171 ); 
   nand2 U3376 ( L6165, L6172, L2823 ); 
   inv U3377 ( L6975, L6981 ); 
   nand2 U3378 ( L6975, L6982, L4058 ); 
   inv U3379 ( L7033, L7039 ); 
   nand2 U3380 ( L7033, L7040, L4063 ); 
   inv U3381 ( L5071, L5077 ); 
   nand2 U3382 ( L5071, L5078, L5080 ); 
   inv U3383 ( L5159, L5165 ); 
   nand2 U3384 ( L5159, L5166, L5090 ); 
   inv U3385 ( L5641, L5647 ); 
   nand2 U3386 ( L5641, L5648, L5650 ); 
   inv U3387 ( L5729, L5735 ); 
   nand2 U3388 ( L5729, L5736, L5660 ); 
   inv U3389 ( L6223, L6229 ); 
   nand2 U3390 ( L6223, L6230, L6232 ); 
   nand2 U3391 ( L6319, L6320, L6321 ); 
   nand2 U3392 ( L7099, L7100, L7101 ); 
   nand2 U3393 ( L7187, L7188, L7189 ); 
   nand2 U3394 ( L6110, L6113, L2817 ); 
   nand2 U3395 ( L6168, L6171, L2822 ); 
   nand2 U3396 ( L6978, L6981, L4057 ); 
   nand2 U3397 ( L7036, L7039, L4062 ); 
   nand2 U3398 ( L5074, L5077, L5079 ); 
   nand2 U3399 ( L5162, L5165, L5089 ); 
   nand2 U3400 ( L5644, L5647, L5649 ); 
   nand2 U3401 ( L5732, L5735, L5659 ); 
   nand2 U3402 ( L6226, L6229, L6231 ); 
   and3 U3403 ( L1762, L1730, L1771, L1782 ); 
   and3 U3404 ( L1757, L1726, L1771, L1783 ); 
   and3 U3405 ( L1762, L1751, L1766, L1784 ); 
   and3 U3406 ( L1757, L1754, L1766, L1785 ); 
   nand2 U3407 ( L2817, L2818, L2819 ); 
   nand2 U3408 ( L2822, L2823, L2824 ); 
   nand2 U3409 ( L4057, L4058, L4059 ); 
   nand2 U3410 ( L4062, L4063, L4064 ); 
   nand2 U3411 ( L5079, L5080, L5081 ); 
   nand2 U3412 ( L5089, L5090, L5091 ); 
   nand2 U3413 ( L5649, L5650, L5651 ); 
   nand2 U3414 ( L5659, L5660, L5661 ); 
   nand2 U3415 ( L6231, L6232, L6233 ); 
   inv U3416 ( L6321, L6327 ); 
   nand2 U3417 ( L6321, L6328, L6252 ); 
   inv U3418 ( L7101, L7107 ); 
   nand2 U3419 ( L7101, L7108, L7110 ); 
   inv U3420 ( L7189, L7195 ); 
   nand2 U3421 ( L7189, L7196, L7120 ); 
   or4 U3422 ( L1782, L1783, L1784, L1785, L5737 ); 
   nand2 U3423 ( L6324, L6327, L6251 ); 
   nand2 U3424 ( L7104, L7107, L7109 ); 
   nand2 U3425 ( L7192, L7195, L7119 ); 
   inv U3426 ( L5081, L5087 ); 
   nand2 U3427 ( L5081, L5088, L985 ); 
   inv U3428 ( L5091, L5097 ); 
   nand2 U3429 ( L5091, L5098, L988 ); 
   inv U3430 ( L5651, L5657 ); 
   nand2 U3431 ( L5651, L5658, L1776 ); 
   inv U3432 ( L5661, L5667 ); 
   nand2 U3433 ( L5661, L5668, L1779 ); 
   and3 U3434 ( L2824, L2784, L2833, L2844 ); 
   and3 U3435 ( L2819, L2780, L2833, L2845 ); 
   and3 U3436 ( L2824, L2813, L2828, L2846 ); 
   and3 U3437 ( L2819, L2816, L2828, L2847 ); 
   and3 U3438 ( L4064, L4032, L4072, L4083 ); 
   and3 U3439 ( L4059, L4028, L4072, L4084 ); 
   and3 U3440 ( L4064, L4053, L4067, L4085 ); 
   and3 U3441 ( L4059, L4056, L4067, L4086 ); 
   inv U3442 ( L6233, L6239 ); 
   nand2 U3443 ( L6233, L6240, L6242 ); 
   nand2 U3444 ( L6251, L6252, L6253 ); 
   nand2 U3445 ( L7109, L7110, L7111 ); 
   nand2 U3446 ( L7119, L7120, L7121 ); 
   nand2 U3447 ( L5084, L5087, L984 ); 
   nand2 U3448 ( L5094, L5097, L987 ); 
   nand2 U3449 ( L5654, L5657, L1775 ); 
   nand2 U3450 ( L5664, L5667, L1778 ); 
   inv U3451 ( L5737, L5743 ); 
   nand2 U3452 ( L6236, L6239, L6241 ); 
   or4 U3453 ( L2844, L2845, L2846, L2847, L6329 ); 
   or4 U3454 ( L4083, L4084, L4085, L4086, L7197 ); 
   nand2 U3455 ( L984, L985, L986 ); 
   nand2 U3456 ( L987, L988, L989 ); 
   nand2 U3457 ( L1775, L1776, L1777 ); 
   nand2 U3458 ( L1778, L1779, L1780 ); 
   inv U3459 ( L6253, L6259 ); 
   nand2 U3460 ( L6253, L6260, L2841 ); 
   inv U3461 ( L7111, L7117 ); 
   nand2 U3462 ( L7111, L7118, L4077 ); 
   inv U3463 ( L7121, L7127 ); 
   nand2 U3464 ( L7121, L7128, L4080 ); 
   nand2 U3465 ( L6241, L6242, L6243 ); 
   inv U3466 ( L989, L990 ); 
   and2 U3467 ( L975, L986, L996 ); 
   inv U3468 ( L1780, L1781 ); 
   and2 U3469 ( L1766, L1777, L1787 ); 
   nand2 U3470 ( L6256, L6259, L2840 ); 
   inv U3471 ( L6329, L6335 ); 
   nand2 U3472 ( L7114, L7117, L4076 ); 
   nand2 U3473 ( L7124, L7127, L4079 ); 
   inv U3474 ( L7197, L7203 ); 
   and2 U3475 ( L990, L980, L995 ); 
   and2 U3476 ( L1781, L1771, L1786 ); 
   inv U3477 ( L6243, L6249 ); 
   nand2 U3478 ( L6243, L6250, L2838 ); 
   nand2 U3479 ( L2840, L2841, L2842 ); 
   nand2 U3480 ( L4076, L4077, L4078 ); 
   nand2 U3481 ( L4079, L4080, L4081 ); 
   nand2 U3482 ( L6246, L6249, L2837 ); 
   inv U3483 ( L2842, L2843 ); 
   inv U3484 ( L4081, L4082 ); 
   and2 U3485 ( L4067, L4078, L4088 ); 
   or2 U3486 ( L995, L996, L5170 ); 
   or2 U3487 ( L1786, L1787, L5740 ); 
   nand2 U3488 ( L2837, L2838, L2839 ); 
   and2 U3489 ( L2843, L2833, L2848 ); 
   and2 U3490 ( L4082, L4072, L4087 ); 
   nand2 U3491 ( L5740, L5743, L1791 ); 
   nand2 U3492 ( L5170, L5173, L1003 ); 
   inv U3493 ( L5170, L5174 ); 
   inv U3494 ( L5740, L5744 ); 
   and2 U3495 ( L2828, L2839, L2849 ); 
   or2 U3496 ( L4087, L4088, L7200 ); 
   nand2 U3497 ( L5737, L5744, L1792 ); 
   nand2 U3498 ( L5167, L5174, L1004 ); 
   or2 U3499 ( L2848, L2849, L6332 ); 
   nand2 U3500 ( L1791, L1792, L320 ); 
   nand2 U3501 ( L1003, L1004, L337 ); 
   nand2 U3502 ( L7200, L7203, L4092 ); 
   inv U3503 ( L7200, L7204 ); 
   inv U3504 ( L320, L321 ); 
   inv U3505 ( L337, L338 ); 
   nand2 U3506 ( L7197, L7204, L4093 ); 
   nand2 U3507 ( L6332, L6335, L2855 ); 
   inv U3508 ( L6332, L6336 ); 
   nand2 U3509 ( L4092, L4093, L369 ); 
   nand2 U3510 ( L6329, L6336, L2856 ); 
   inv U3511 ( L369, L370 ); 
   nand2 U3512 ( L2855, L2856, L398 ); 
   inv U3513 ( L398, L399 ); 
endmodule

