/****************************************************************************
 *                                                                          *
 *  VERILOG VERSION of ORIGINAL NETLIST for c3540                           *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *                                                                          *
 *                Sep 16, 1998                                              *
 *                                                                          *
****************************************************************************/

module c3540g (
        L50, L58, L68, L77, L87, L97, L107,
        L116, L226, L232, L238, L244, L250, L257, L264,
        L270, L124, L125, L128, L132, L137, L143, L150,
        L159, L283, L294, L303, L311, L317, L322, L326,
        L329, L222, L223, L330, L274, L2897, L200, L190,
        L179, L343, L213, L169, L45, L41, L1698, L33,
        L20, L13, L1,
        L375, L378, L381, L384, L387, L390, L393,
        L396, L407, L409, L402, L351, L358, L405, L399,
        L369, L372, L353, L355, L361, L364, L367);
 
   input
        L50, L58, L68, L77, L87, L97, L107,
        L116, L226, L232, L238, L244, L250, L257, L264,
        L270, L124, L125, L128, L132, L137, L143, L150,
        L159, L283, L294, L303, L311, L317, L322, L326,
        L329, L222, L223, L330, L274, L2897, L200, L190,
        L179, L343, L213, L169, L45, L41, L1698, L33,
        L20, L13, L1;
 
   output
        L375, L378, L381, L384, L387, L390, L393,
        L396, L407, L409, L402, L351, L358, L405, L399,
        L369, L372, L353, L355, L361, L364, L367;



   buffer U1 ( L50, L432 ); 
   inv U2 ( L50, L442 ); 
   buffer U3 ( L58, L447 ); 
   inv U4 ( L58, L456 ); 
   buffer U5 ( L68, L460 ); 
   inv U6 ( L68, L463 ); 
   buffer U7 ( L68, L467 ); 
   buffer U8 ( L77, L476 ); 
   inv U9 ( L77, L479 ); 
   buffer U10 ( L77, L483 ); 
   buffer U11 ( L87, L492 ); 
   inv U12 ( L87, L501 ); 
   buffer U13 ( L97, L504 ); 
   inv U14 ( L97, L513 ); 
   buffer U15 ( L107, L517 ); 
   inv U16 ( L107, L526 ); 
   buffer U17 ( L116, L530 ); 
   inv U18 ( L116, L540 ); 
   or2 U19 ( L257, L264, L587 ); 
   inv U20 ( L1, L704 ); 
   buffer U21 ( L1, L707 ); 
   inv U22 ( L1, L714 ); 
   buffer U23 ( L13, L717 ); 
   inv U24 ( L13, L724 ); 
   and2 U25 ( L13, L20, L731 ); 
   inv U26 ( L20, L732 ); 
   buffer U27 ( L20, L736 ); 
   inv U28 ( L20, L741 ); 
   inv U29 ( L33, L758 ); 
   buffer U30 ( L33, L776 ); 
   inv U31 ( L33, L780 ); 
   and2 U32 ( L33, L41, L788 ); 
   inv U33 ( L41, L791 ); 
   or2 U34 ( L41, L45, L798 ); 
   buffer U35 ( L45, L799 ); 
   inv U36 ( L45, L802 ); 
   inv U37 ( L50, L826 ); 
   buffer U38 ( L58, L828 ); 
   inv U39 ( L58, L831 ); 
   buffer U40 ( L68, L833 ); 
   inv U41 ( L68, L836 ); 
   buffer U42 ( L87, L839 ); 
   inv U43 ( L87, L842 ); 
   buffer U44 ( L97, L845 ); 
   inv U45 ( L97, L848 ); 
   inv U46 ( L107, L851 ); 
   buffer U47 ( L1, L890 ); 
   buffer U48 ( L68, L898 ); 
   buffer U49 ( L107, L907 ); 
   inv U50 ( L20, L1032 ); 
   buffer U51 ( L190, L1035 ); 
   inv U52 ( L200, L1048 ); 
   and2 U53 ( L20, L200, L1049 ); 
   nand2 U54 ( L20, L200, L1050 ); 
   and2 U55 ( L20, L179, L1051 ); 
   inv U56 ( L20, L1540 ); 
   or2 U57 ( L1698, L33, L1699 ); 
   nand2 U58 ( L1, L13, L1826 ); 
   nand3 U59 ( L1, L20, L33, L1827 ); 
   inv U60 ( L20, L1828 ); 
   inv U61 ( L33, L2051 ); 
   buffer U62 ( L179, L2478 ); 
   inv U63 ( L213, L2865 ); 
   buffer U64 ( L343, L2868 ); 
   buffer U65 ( L226, L2931 ); 
   buffer U66 ( L232, L2934 ); 
   buffer U67 ( L238, L2939 ); 
   buffer U68 ( L244, L2942 ); 
   buffer U69 ( L250, L2947 ); 
   buffer U70 ( L257, L2950 ); 
   buffer U71 ( L264, L2957 ); 
   buffer U72 ( L270, L2960 ); 
   buffer U73 ( L50, L3007 ); 
   buffer U74 ( L58, L3079 ); 
   buffer U75 ( L58, L3087 ); 
   buffer U76 ( L97, L3095 ); 
   buffer U77 ( L97, L3103 ); 
   buffer U78 ( L330, L3419 ); 
   and2 U79 ( L250, L587, L588 ); 
   or2 U80 ( L758, L20, L759 ); 
   or2 U81 ( L1540, L169, L1541 ); 
   inv U82 ( L731, L1772 ); 
   or2 U83 ( L1828, L1, L1829 ); 
   and2 U84 ( L1826, L1827, L1834 ); 
   or2 U85 ( L2051, L1, L2052 ); 
   and3 U86 ( L826, L831, L836, L625 ); 
   nand2 U87 ( L226, L432, L545 ); 
   nand2 U88 ( L232, L447, L546 ); 
   nand2 U89 ( L238, L467, L547 ); 
   nand2 U90 ( L244, L483, L548 ); 
   nand2 U91 ( L250, L492, L549 ); 
   nand2 U92 ( L257, L504, L550 ); 
   nand2 U93 ( L264, L517, L551 ); 
   nand2 U94 ( L270, L530, L552 ); 
   inv U95 ( L2931, L2937 ); 
   inv U96 ( L2934, L2938 ); 
   inv U97 ( L2939, L2945 ); 
   inv U98 ( L2942, L2946 ); 
   nand2 U99 ( L456, L463, L621 ); 
   nand2 U100 ( L513, L526, L626 ); 
   nand2 U101 ( L460, L476, L635 ); 
   buffer U102 ( L442, L636 ); 
   inv U103 ( L3079, L3085 ); 
   inv U104 ( L3095, L3101 ); 
   buffer U105 ( L802, L657 ); 
   buffer U106 ( L802, L675 ); 
   buffer U107 ( L717, L721 ); 
   buffer U108 ( L780, L784 ); 
   buffer U109 ( L791, L794 ); 
   and2 U110 ( L714, L798, L807 ); 
   and3 U111 ( L714, L799, L791, L816 ); 
   and2 U112 ( L704, L799, L823 ); 
   and3 U113 ( L707, L724, L736, L860 ); 
   nand3 U114 ( L707, L724, L736, L861 ); 
   nand2 U115 ( L707, L724, L864 ); 
   buffer U116 ( L890, L893 ); 
   nand3 U117 ( L717, L732, L45, L896 ); 
   nand3 U118 ( L826, L831, L836, L897 ); 
   inv U119 ( L3087, L3093 ); 
   and3 U120 ( L842, L848, L851, L905 ); 
   nand3 U121 ( L842, L848, L851, L906 ); 
   inv U122 ( L3103, L3109 ); 
   inv U123 ( L741, L973 ); 
   inv U124 ( L741, L980 ); 
   inv U125 ( L741, L987 ); 
   inv U126 ( L741, L994 ); 
   inv U127 ( L741, L1001 ); 
   inv U128 ( L741, L1008 ); 
   inv U129 ( L741, L1015 ); 
   inv U130 ( L741, L1022 ); 
   or2 U131 ( L1032, L1035, L1038 ); 
   nor2 U132 ( L1032, L1035, L1043 ); 
   buffer U133 ( L1051, L1054 ); 
   inv U134 ( L1051, L1057 ); 
   buffer U135 ( L776, L1512 ); 
   buffer U136 ( L780, L1681 ); 
   inv U137 ( L1699, L1717 ); 
   inv U138 ( L1699, L1724 ); 
   inv U139 ( L1699, L1731 ); 
   inv U140 ( L1699, L1738 ); 
   inv U141 ( L1699, L1745 ); 
   inv U142 ( L1699, L1752 ); 
   inv U143 ( L1699, L1759 ); 
   inv U144 ( L1699, L1766 ); 
   or2 U145 ( L1, L1772, L1773 ); 
   inv U146 ( L788, L1790 ); 
   inv U147 ( L788, L1808 ); 
   and3 U148 ( L704, L717, L732, L2278 ); 
   inv U149 ( L2478, L2481 ); 
   inv U150 ( L3419, L3425 ); 
   or2 U151 ( L2865, L2868, L2871 ); 
   nor2 U152 ( L2865, L2868, L2874 ); 
   inv U153 ( L2947, L2953 ); 
   inv U154 ( L2950, L2954 ); 
   inv U155 ( L2957, L2963 ); 
   inv U156 ( L2960, L2964 ); 
   buffer U157 ( L456, L3010 ); 
   inv U158 ( L3007, L3013 ); 
   buffer U159 ( L463, L3017 ); 
   buffer U160 ( L479, L3020 ); 
   buffer U161 ( L501, L3027 ); 
   buffer U162 ( L513, L3030 ); 
   buffer U163 ( L526, L3037 ); 
   buffer U164 ( L540, L3040 ); 
   buffer U165 ( L898, L3082 ); 
   buffer U166 ( L898, L3090 ); 
   buffer U167 ( L907, L3098 ); 
   buffer U168 ( L907, L3106 ); 
   nand2 U169 ( L479, L625, L352 ); 
   and4 U170 ( L545, L546, L547, L548, L553 ); 
   and4 U171 ( L549, L550, L551, L552, L554 ); 
   nand2 U172 ( L2934, L2937, L555 ); 
   nand2 U173 ( L2931, L2938, L556 ); 
   nand2 U174 ( L2942, L2945, L560 ); 
   nand2 U175 ( L2939, L2946, L561 ); 
   and2 U176 ( L432, L621, L650 ); 
   and2 U177 ( L890, L896, L956 ); 
   inv U178 ( L759, L974 ); 
   and2 U179 ( L741, L759, L975 ); 
   and2 U180 ( L897, L973, L976 ); 
   inv U181 ( L759, L981 ); 
   and2 U182 ( L741, L759, L982 ); 
   inv U183 ( L759, L988 ); 
   and2 U184 ( L741, L759, L989 ); 
   and2 U185 ( L836, L987, L990 ); 
   inv U186 ( L759, L995 ); 
   and2 U187 ( L741, L759, L996 ); 
   and2 U188 ( L77, L994, L997 ); 
   inv U189 ( L759, L1002 ); 
   and2 U190 ( L741, L759, L1003 ); 
   and2 U191 ( L906, L1001, L1004 ); 
   inv U192 ( L759, L1009 ); 
   and2 U193 ( L741, L759, L1010 ); 
   inv U194 ( L759, L1016 ); 
   and2 U195 ( L741, L759, L1017 ); 
   and2 U196 ( L851, L1015, L1018 ); 
   inv U197 ( L759, L1023 ); 
   and2 U198 ( L741, L759, L1024 ); 
   and2 U199 ( L116, L1022, L1025 ); 
   and2 U200 ( L222, L1717, L1720 ); 
   and2 U201 ( L223, L1724, L1727 ); 
   and2 U202 ( L226, L1731, L1734 ); 
   and2 U203 ( L232, L1738, L1741 ); 
   and2 U204 ( L238, L1745, L1748 ); 
   and2 U205 ( L244, L1752, L1755 ); 
   and2 U206 ( L250, L1759, L1762 ); 
   and2 U207 ( L257, L1766, L1769 ); 
   and3 U208 ( L1, L13, L1790, L1791 ); 
   and3 U209 ( L1, L13, L1808, L1809 ); 
   inv U210 ( L1834, L1851 ); 
   inv U211 ( L1834, L1901 ); 
   inv U212 ( L1834, L1952 ); 
   inv U213 ( L1834, L2002 ); 
   inv U214 ( L1834, L2057 ); 
   inv U215 ( L1834, L2109 ); 
   inv U216 ( L1834, L2162 ); 
   inv U217 ( L1834, L2214 ); 
   nand2 U218 ( L2950, L2953, L2955 ); 
   nand2 U219 ( L2947, L2954, L2956 ); 
   nand2 U220 ( L2960, L2963, L2965 ); 
   nand2 U221 ( L2957, L2964, L2966 ); 
   inv U222 ( L352, L353 ); 
   and2 U223 ( L87, L626, L354 ); 
   nand2 U224 ( L555, L556, L557 ); 
   nand2 U225 ( L560, L561, L562 ); 
   nand2 U226 ( L553, L554, L586 ); 
   and2 U227 ( L540, L905, L630 ); 
   nand2 U228 ( L540, L905, L634 ); 
   inv U229 ( L636, L639 ); 
   nand2 U230 ( L3082, L3085, L642 ); 
   inv U231 ( L3082, L3086 ); 
   and2 U232 ( L460, L636, L644 ); 
   nand2 U233 ( L3098, L3101, L646 ); 
   inv U234 ( L3098, L3102 ); 
   nand2 U235 ( L87, L626, L654 ); 
   inv U236 ( L657, L660 ); 
   inv U237 ( L675, L678 ); 
   nand2 U238 ( L860, L776, L804 ); 
   nand2 U239 ( L860, L780, L806 ); 
   nand3 U240 ( L707, L721, L736, L855 ); 
   nand4 U241 ( L707, L724, L736, L794, L867 ); 
   nand2 U242 ( L3090, L3093, L903 ); 
   inv U243 ( L3090, L3094 ); 
   nand2 U244 ( L3106, L3109, L912 ); 
   inv U245 ( L3106, L3110 ); 
   inv U246 ( L861, L915 ); 
   inv U247 ( L893, L927 ); 
   inv U248 ( L864, L941 ); 
   and2 U249 ( L828, L974, L977 ); 
   and2 U250 ( L150, L975, L978 ); 
   and2 U251 ( L833, L981, L984 ); 
   and2 U252 ( L159, L982, L985 ); 
   and2 U253 ( L77, L988, L991 ); 
   and2 U254 ( L50, L989, L992 ); 
   and2 U255 ( L839, L995, L998 ); 
   and2 U256 ( L828, L996, L999 ); 
   and2 U257 ( L845, L1002, L1005 ); 
   and2 U258 ( L833, L1003, L1006 ); 
   and2 U259 ( L107, L1009, L1012 ); 
   and2 U260 ( L77, L1010, L1013 ); 
   and2 U261 ( L116, L1016, L1019 ); 
   and2 U262 ( L839, L1017, L1020 ); 
   and2 U263 ( L283, L1023, L1026 ); 
   and2 U264 ( L845, L1024, L1027 ); 
   and2 U265 ( L200, L1054, L1060 ); 
   and2 U266 ( L1048, L1054, L1063 ); 
   and2 U267 ( L1049, L1057, L1066 ); 
   and2 U268 ( L1050, L1057, L1069 ); 
   nand2 U269 ( L784, L794, L1527 ); 
   nand2 U270 ( L776, L794, L1530 ); 
   nand3 U271 ( L707, L721, L1541, L1542 ); 
   nand3 U272 ( L724, L732, L784, L1563 ); 
   nand2 U273 ( L724, L784, L1572 ); 
   inv U274 ( L1512, L1581 ); 
   inv U275 ( L1512, L1585 ); 
   inv U276 ( L1512, L1589 ); 
   inv U277 ( L1512, L1593 ); 
   inv U278 ( L1512, L1597 ); 
   inv U279 ( L1512, L1601 ); 
   inv U280 ( L1512, L1605 ); 
   inv U281 ( L1681, L1716 ); 
   and2 U282 ( L1681, L1699, L1718 ); 
   inv U283 ( L1681, L1723 ); 
   and2 U284 ( L1681, L1699, L1725 ); 
   inv U285 ( L1681, L1730 ); 
   and2 U286 ( L1681, L1699, L1732 ); 
   inv U287 ( L1681, L1737 ); 
   and2 U288 ( L1681, L1699, L1739 ); 
   inv U289 ( L1681, L1744 ); 
   and2 U290 ( L1681, L1699, L1746 ); 
   inv U291 ( L1681, L1751 ); 
   and2 U292 ( L1681, L1699, L1753 ); 
   inv U293 ( L1681, L1758 ); 
   and2 U294 ( L1681, L1699, L1760 ); 
   inv U295 ( L1681, L1765 ); 
   and2 U296 ( L1681, L1699, L1767 ); 
   and2 U297 ( L1834, L1773, L1852 ); 
   nor2 U298 ( L50, L1773, L1856 ); 
   inv U299 ( L807, L1870 ); 
   and2 U300 ( L1834, L1773, L1902 ); 
   nor2 U301 ( L58, L1773, L1906 ); 
   inv U302 ( L807, L1920 ); 
   and2 U303 ( L1834, L1773, L1953 ); 
   nor2 U304 ( L68, L1773, L1957 ); 
   inv U305 ( L807, L1971 ); 
   and2 U306 ( L1834, L1773, L2003 ); 
   nor2 U307 ( L77, L1773, L2007 ); 
   inv U308 ( L807, L2021 ); 
   and2 U309 ( L1834, L1773, L2058 ); 
   nor2 U310 ( L87, L1773, L2062 ); 
   inv U311 ( L823, L2076 ); 
   and2 U312 ( L1834, L1773, L2110 ); 
   nor2 U313 ( L97, L1773, L2114 ); 
   inv U314 ( L816, L2128 ); 
   and2 U315 ( L1834, L1773, L2163 ); 
   nor2 U316 ( L107, L1773, L2167 ); 
   inv U317 ( L816, L2181 ); 
   and2 U318 ( L1834, L1773, L2215 ); 
   nor2 U319 ( L116, L1773, L2219 ); 
   inv U320 ( L816, L2233 ); 
   and2 U321 ( L2278, L213, L2285 ); 
   nand2 U322 ( L2278, L213, L2288 ); 
   and3 U323 ( L2278, L213, L343, L2289 ); 
   nand3 U324 ( L2278, L213, L343, L2293 ); 
   and3 U325 ( L2278, L213, L343, L2298 ); 
   nand3 U326 ( L2278, L213, L343, L2302 ); 
   buffer U327 ( L2874, L2877 ); 
   nand2 U328 ( L2955, L2956, L2983 ); 
   nand2 U329 ( L2965, L2966, L2986 ); 
   inv U330 ( L3010, L3014 ); 
   nand2 U331 ( L3010, L3013, L3015 ); 
   inv U332 ( L3017, L3023 ); 
   inv U333 ( L3020, L3024 ); 
   inv U334 ( L3027, L3033 ); 
   inv U335 ( L3030, L3034 ); 
   inv U336 ( L3037, L3043 ); 
   inv U337 ( L3040, L3044 ); 
   inv U338 ( L354, L355 ); 
   nand2 U339 ( L3079, L3086, L643 ); 
   nand2 U340 ( L3095, L3102, L647 ); 
   and2 U341 ( L650, L675, L680 ); 
   nand2 U342 ( L3087, L3094, L904 ); 
   nand2 U343 ( L3103, L3110, L913 ); 
   and2 U344 ( L588, L915, L920 ); 
   or3 U345 ( L976, L977, L978, L979 ); 
   or3 U346 ( L990, L991, L992, L993 ); 
   or3 U347 ( L997, L998, L999, L1000 ); 
   or3 U348 ( L1004, L1005, L1006, L1007 ); 
   or3 U349 ( L1018, L1019, L1020, L1021 ); 
   or3 U350 ( L1025, L1026, L1027, L1028 ); 
   and2 U351 ( L77, L1716, L1719 ); 
   and2 U352 ( L223, L1718, L1721 ); 
   and2 U353 ( L87, L1723, L1726 ); 
   and2 U354 ( L226, L1725, L1728 ); 
   and2 U355 ( L97, L1730, L1733 ); 
   and2 U356 ( L232, L1732, L1735 ); 
   and2 U357 ( L107, L1737, L1740 ); 
   and2 U358 ( L238, L1739, L1742 ); 
   and2 U359 ( L116, L1744, L1747 ); 
   and2 U360 ( L244, L1746, L1749 ); 
   and2 U361 ( L283, L1751, L1754 ); 
   and2 U362 ( L250, L1753, L1756 ); 
   and2 U363 ( L294, L1758, L1761 ); 
   and2 U364 ( L257, L1760, L1763 ); 
   and2 U365 ( L303, L1765, L1768 ); 
   and2 U366 ( L264, L1767, L1770 ); 
   buffer U367 ( L1791, L1794 ); 
   inv U368 ( L1791, L1799 ); 
   buffer U369 ( L1809, L1812 ); 
   inv U370 ( L1809, L1817 ); 
   and3 U371 ( L50, L1829, L1852, L1859 ); 
   and3 U372 ( L58, L1829, L1902, L1909 ); 
   and3 U373 ( L68, L1829, L1953, L1960 ); 
   and3 U374 ( L77, L1829, L2003, L2010 ); 
   and3 U375 ( L87, L2052, L2058, L2065 ); 
   and3 U376 ( L97, L2052, L2110, L2117 ); 
   and3 U377 ( L107, L2052, L2163, L2170 ); 
   and3 U378 ( L116, L2052, L2215, L2222 ); 
   inv U379 ( L956, L2678 ); 
   inv U380 ( L956, L2697 ); 
   inv U381 ( L956, L2716 ); 
   inv U382 ( L956, L2733 ); 
   inv U383 ( L956, L2751 ); 
   inv U384 ( L956, L2768 ); 
   inv U385 ( L956, L2785 ); 
   inv U386 ( L956, L2802 ); 
   nand2 U387 ( L3007, L3014, L3016 ); 
   nand2 U388 ( L3020, L3023, L3025 ); 
   nand2 U389 ( L3017, L3024, L3026 ); 
   nand2 U390 ( L3030, L3033, L3035 ); 
   nand2 U391 ( L3027, L3034, L3036 ); 
   nand2 U392 ( L3040, L3043, L3045 ); 
   nand2 U393 ( L3037, L3044, L3046 ); 
   inv U394 ( L2983, L2989 ); 
   inv U395 ( L2986, L2990 ); 
   inv U396 ( L804, L610 ); 
   and2 U397 ( L804, L806, L613 ); 
   inv U398 ( L806, L616 ); 
   nand2 U399 ( L642, L643, L640 ); 
   nand2 U400 ( L646, L647, L648 ); 
   and4 U401 ( L630, L635, L442, L58, L655 ); 
   inv U402 ( L804, L665 ); 
   and2 U403 ( L804, L806, L668 ); 
   inv U404 ( L806, L671 ); 
   inv U405 ( L804, L683 ); 
   inv U406 ( L806, L685 ); 
   and2 U407 ( L804, L806, L688 ); 
   inv U408 ( L804, L694 ); 
   inv U409 ( L806, L696 ); 
   and2 U410 ( L804, L806, L699 ); 
   buffer U411 ( L867, L870 ); 
   buffer U412 ( L867, L887 ); 
   nand2 U413 ( L903, L904, L901 ); 
   nand2 U414 ( L912, L913, L910 ); 
   inv U415 ( L855, L914 ); 
   and2 U416 ( L855, L861, L916 ); 
   inv U417 ( L855, L942 ); 
   and2 U418 ( L864, L855, L943 ); 
   nand2 U419 ( L1043, L1069, L1072 ); 
   nand2 U420 ( L1043, L1066, L1084 ); 
   nand2 U421 ( L1038, L1069, L1096 ); 
   nand2 U422 ( L1038, L1066, L1108 ); 
   nand2 U423 ( L1043, L1063, L1120 ); 
   nand2 U424 ( L1043, L1060, L1132 ); 
   nand2 U425 ( L1038, L1063, L1144 ); 
   nand2 U426 ( L1038, L1060, L1156 ); 
   inv U427 ( L1527, L1533 ); 
   inv U428 ( L1530, L1534 ); 
   and2 U429 ( L1527, L1530, L1535 ); 
   buffer U430 ( L1542, L1545 ); 
   buffer U431 ( L1542, L1554 ); 
   inv U432 ( L1572, L1610 ); 
   inv U433 ( L1572, L1619 ); 
   inv U434 ( L1572, L1628 ); 
   inv U435 ( L1572, L1637 ); 
   inv U436 ( L1563, L1646 ); 
   inv U437 ( L1563, L1655 ); 
   inv U438 ( L1563, L1664 ); 
   inv U439 ( L1563, L1673 ); 
   or3 U440 ( L1719, L1720, L1721, L1722 ); 
   or3 U441 ( L1726, L1727, L1728, L1729 ); 
   or3 U442 ( L1733, L1734, L1735, L1736 ); 
   or3 U443 ( L1740, L1741, L1742, L1743 ); 
   or3 U444 ( L1747, L1748, L1749, L1750 ); 
   or3 U445 ( L1754, L1755, L1756, L1757 ); 
   or3 U446 ( L1761, L1762, L1763, L1764 ); 
   or3 U447 ( L1768, L1769, L1770, L1771 ); 
   and2 U448 ( L979, L1851, L1853 ); 
   and2 U449 ( L993, L1952, L1954 ); 
   and2 U450 ( L1000, L2002, L2004 ); 
   and2 U451 ( L1007, L2057, L2059 ); 
   and2 U452 ( L1021, L2162, L2164 ); 
   and2 U453 ( L1028, L2214, L2216 ); 
   buffer U454 ( L2293, L2485 ); 
   and2 U455 ( L2877, L2897, L2900 ); 
   nand2 U456 ( L2877, L2897, L2903 ); 
   buffer U457 ( L557, L2967 ); 
   buffer U458 ( L562, L2970 ); 
   buffer U459 ( L557, L2975 ); 
   buffer U460 ( L562, L2978 ); 
   nand2 U461 ( L3015, L3016, L3047 ); 
   nand2 U462 ( L3025, L3026, L3050 ); 
   nand2 U463 ( L3035, L3036, L3055 ); 
   nand2 U464 ( L3045, L3046, L3058 ); 
   nand2 U465 ( L2986, L2989, L574 ); 
   nand2 U466 ( L2983, L2990, L575 ); 
   and2 U467 ( L501, L613, L617 ); 
   and3 U468 ( L640, L476, L639, L641 ); 
   and2 U469 ( L530, L648, L649 ); 
   and2 U470 ( L655, L657, L662 ); 
   and2 U471 ( L513, L668, L672 ); 
   and2 U472 ( L654, L685, L690 ); 
   and2 U473 ( L540, L688, L691 ); 
   and2 U474 ( L634, L696, L701 ); 
   and2 U475 ( L526, L699, L702 ); 
   inv U476 ( L901, L902 ); 
   inv U477 ( L910, L911 ); 
   and2 U478 ( L650, L914, L917 ); 
   and2 U479 ( L586, L916, L923 ); 
   and2 U480 ( L442, L1535, L1538 ); 
   and3 U481 ( L1817, L226, L1870, L1871 ); 
   and3 U482 ( L1817, L274, L807, L1872 ); 
   and2 U483 ( L1812, L1722, L1873 ); 
   and3 U484 ( L1817, L232, L1920, L1921 ); 
   and3 U485 ( L1817, L274, L807, L1922 ); 
   and2 U486 ( L1812, L1729, L1923 ); 
   and3 U487 ( L1817, L238, L1971, L1972 ); 
   and3 U488 ( L1817, L274, L807, L1973 ); 
   and2 U489 ( L1812, L1736, L1974 ); 
   and3 U490 ( L1817, L244, L2021, L2022 ); 
   and3 U491 ( L1817, L274, L807, L2023 ); 
   and2 U492 ( L1812, L1743, L2024 ); 
   and3 U493 ( L1799, L250, L2076, L2077 ); 
   and3 U494 ( L1799, L274, L823, L2078 ); 
   and2 U495 ( L1794, L1750, L2079 ); 
   and3 U496 ( L1799, L257, L2128, L2129 ); 
   and3 U497 ( L1799, L274, L816, L2130 ); 
   and2 U498 ( L1794, L1757, L2131 ); 
   and3 U499 ( L1799, L264, L2181, L2182 ); 
   and3 U500 ( L1799, L274, L816, L2183 ); 
   and2 U501 ( L1794, L1764, L2184 ); 
   and3 U502 ( L1799, L270, L2233, L2234 ); 
   and3 U503 ( L1799, L274, L816, L2235 ); 
   and2 U504 ( L1794, L1771, L2236 ); 
   inv U505 ( L2967, L2973 ); 
   inv U506 ( L2970, L2974 ); 
   inv U507 ( L2975, L2981 ); 
   inv U508 ( L2978, L2982 ); 
   nand2 U509 ( L574, L575, L576 ); 
   inv U510 ( L3047, L3053 ); 
   inv U511 ( L3050, L3054 ); 
   inv U512 ( L3055, L3061 ); 
   inv U513 ( L3058, L3062 ); 
   or2 U514 ( L641, L644, L645 ); 
   inv U515 ( L887, L926 ); 
   and2 U516 ( L887, L893, L928 ); 
   and2 U517 ( L649, L942, L947 ); 
   and2 U518 ( L902, L980, L983 ); 
   and2 U519 ( L911, L1008, L1011 ); 
   buffer U520 ( L1072, L1075 ); 
   buffer U521 ( L1084, L1087 ); 
   buffer U522 ( L1096, L1099 ); 
   buffer U523 ( L1108, L1111 ); 
   buffer U524 ( L1120, L1123 ); 
   buffer U525 ( L1132, L1135 ); 
   buffer U526 ( L1144, L1147 ); 
   buffer U527 ( L1156, L1159 ); 
   buffer U528 ( L1072, L1168 ); 
   buffer U529 ( L1084, L1177 ); 
   buffer U530 ( L1096, L1186 ); 
   buffer U531 ( L1108, L1195 ); 
   buffer U532 ( L1120, L1204 ); 
   buffer U533 ( L1132, L1213 ); 
   buffer U534 ( L1144, L1222 ); 
   buffer U535 ( L1156, L1231 ); 
   inv U536 ( L1545, L1609 ); 
   and2 U537 ( L1545, L1572, L1611 ); 
   inv U538 ( L1545, L1618 ); 
   and2 U539 ( L1545, L1572, L1620 ); 
   inv U540 ( L1545, L1627 ); 
   and2 U541 ( L1545, L1572, L1629 ); 
   inv U542 ( L1545, L1636 ); 
   and2 U543 ( L1545, L1572, L1638 ); 
   inv U544 ( L1554, L1645 ); 
   and2 U545 ( L1554, L1563, L1647 ); 
   inv U546 ( L1554, L1654 ); 
   and2 U547 ( L1554, L1563, L1656 ); 
   inv U548 ( L1554, L1663 ); 
   and2 U549 ( L1554, L1563, L1665 ); 
   inv U550 ( L1554, L1672 ); 
   and2 U551 ( L1554, L1563, L1674 ); 
   or3 U552 ( L1853, L1856, L1859, L1862 ); 
   nor3 U553 ( L1853, L1856, L1859, L1866 ); 
   or3 U554 ( L1871, L1872, L1873, L1874 ); 
   or3 U555 ( L1921, L1922, L1923, L1924 ); 
   or3 U556 ( L1954, L1957, L1960, L1963 ); 
   nor3 U557 ( L1954, L1957, L1960, L1967 ); 
   or3 U558 ( L1972, L1973, L1974, L1975 ); 
   or3 U559 ( L2004, L2007, L2010, L2013 ); 
   nor3 U560 ( L2004, L2007, L2010, L2017 ); 
   or3 U561 ( L2022, L2023, L2024, L2025 ); 
   or3 U562 ( L2059, L2062, L2065, L2068 ); 
   nor3 U563 ( L2059, L2062, L2065, L2072 ); 
   or3 U564 ( L2077, L2078, L2079, L2080 ); 
   or3 U565 ( L2129, L2130, L2131, L2132 ); 
   or3 U566 ( L2164, L2167, L2170, L2173 ); 
   nor3 U567 ( L2164, L2167, L2170, L2177 ); 
   or3 U568 ( L2182, L2183, L2184, L2185 ); 
   or3 U569 ( L2216, L2219, L2222, L2225 ); 
   nor3 U570 ( L2216, L2219, L2222, L2229 ); 
   or3 U571 ( L2234, L2235, L2236, L2237 ); 
   inv U572 ( L2485, L2488 ); 
   inv U573 ( L870, L2679 ); 
   and2 U574 ( L956, L870, L2680 ); 
   inv U575 ( L870, L2698 ); 
   and2 U576 ( L956, L870, L2699 ); 
   inv U577 ( L870, L2717 ); 
   and2 U578 ( L956, L870, L2718 ); 
   inv U579 ( L870, L2734 ); 
   and2 U580 ( L956, L870, L2735 ); 
   inv U581 ( L870, L2752 ); 
   and2 U582 ( L956, L870, L2753 ); 
   inv U583 ( L870, L2769 ); 
   and2 U584 ( L956, L870, L2770 ); 
   inv U585 ( L870, L2786 ); 
   and2 U586 ( L956, L870, L2787 ); 
   inv U587 ( L870, L2803 ); 
   and2 U588 ( L956, L870, L2804 ); 
   or3 U589 ( L917, L920, L923, L359 ); 
   nor3 U590 ( L917, L920, L923, L1029 ); 
   nand2 U591 ( L2970, L2973, L565 ); 
   nand2 U592 ( L2967, L2974, L566 ); 
   nand2 U593 ( L2978, L2981, L569 ); 
   nand2 U594 ( L2975, L2982, L570 ); 
   nand2 U595 ( L3050, L3053, L589 ); 
   nand2 U596 ( L3047, L3054, L590 ); 
   nand2 U597 ( L3058, L3061, L595 ); 
   nand2 U598 ( L3055, L3062, L596 ); 
   and2 U599 ( L650, L926, L929 ); 
   and2 U600 ( L630, L928, L938 ); 
   and2 U601 ( L645, L941, L944 ); 
   or3 U602 ( L983, L984, L985, L986 ); 
   or3 U603 ( L1011, L1012, L1013, L1014 ); 
   and2 U604 ( L442, L1611, L1616 ); 
   and2 U605 ( L456, L1620, L1625 ); 
   and2 U606 ( L463, L1629, L1634 ); 
   and2 U607 ( L479, L1638, L1643 ); 
   inv U608 ( L1029, L360 ); 
   nand2 U609 ( L565, L566, L567 ); 
   nand2 U610 ( L569, L570, L571 ); 
   buffer U611 ( L576, L579 ); 
   nand2 U612 ( L589, L590, L591 ); 
   nand2 U613 ( L595, L596, L597 ); 
   and2 U614 ( L576, L610, L614 ); 
   inv U615 ( L1075, L1240 ); 
   inv U616 ( L1087, L1241 ); 
   inv U617 ( L1099, L1242 ); 
   inv U618 ( L1111, L1243 ); 
   inv U619 ( L1123, L1244 ); 
   inv U620 ( L1135, L1245 ); 
   inv U621 ( L1147, L1246 ); 
   inv U622 ( L1159, L1247 ); 
   inv U623 ( L1075, L1257 ); 
   inv U624 ( L1087, L1258 ); 
   inv U625 ( L1099, L1259 ); 
   inv U626 ( L1111, L1260 ); 
   inv U627 ( L1123, L1261 ); 
   inv U628 ( L1135, L1262 ); 
   inv U629 ( L1147, L1263 ); 
   inv U630 ( L1159, L1264 ); 
   inv U631 ( L1075, L1274 ); 
   inv U632 ( L1087, L1275 ); 
   inv U633 ( L1099, L1276 ); 
   inv U634 ( L1111, L1277 ); 
   inv U635 ( L1123, L1278 ); 
   inv U636 ( L1135, L1279 ); 
   inv U637 ( L1147, L1280 ); 
   inv U638 ( L1159, L1281 ); 
   inv U639 ( L1075, L1291 ); 
   inv U640 ( L1087, L1292 ); 
   inv U641 ( L1099, L1293 ); 
   inv U642 ( L1111, L1294 ); 
   inv U643 ( L1123, L1295 ); 
   inv U644 ( L1135, L1296 ); 
   inv U645 ( L1147, L1297 ); 
   inv U646 ( L1159, L1298 ); 
   inv U647 ( L1075, L1308 ); 
   inv U648 ( L1087, L1309 ); 
   inv U649 ( L1099, L1310 ); 
   inv U650 ( L1111, L1311 ); 
   inv U651 ( L1123, L1312 ); 
   inv U652 ( L1135, L1313 ); 
   inv U653 ( L1147, L1314 ); 
   inv U654 ( L1159, L1315 ); 
   inv U655 ( L1075, L1325 ); 
   inv U656 ( L1087, L1326 ); 
   inv U657 ( L1099, L1327 ); 
   inv U658 ( L1111, L1328 ); 
   inv U659 ( L1123, L1329 ); 
   inv U660 ( L1135, L1330 ); 
   inv U661 ( L1147, L1331 ); 
   inv U662 ( L1159, L1332 ); 
   inv U663 ( L1075, L1342 ); 
   inv U664 ( L1087, L1343 ); 
   inv U665 ( L1099, L1344 ); 
   inv U666 ( L1111, L1345 ); 
   inv U667 ( L1123, L1346 ); 
   inv U668 ( L1135, L1347 ); 
   inv U669 ( L1147, L1348 ); 
   inv U670 ( L1159, L1349 ); 
   inv U671 ( L1075, L1359 ); 
   inv U672 ( L1087, L1360 ); 
   inv U673 ( L1099, L1361 ); 
   inv U674 ( L1111, L1362 ); 
   inv U675 ( L1123, L1363 ); 
   inv U676 ( L1135, L1364 ); 
   inv U677 ( L1147, L1365 ); 
   inv U678 ( L1159, L1366 ); 
   inv U679 ( L1168, L1376 ); 
   inv U680 ( L1177, L1377 ); 
   inv U681 ( L1186, L1378 ); 
   inv U682 ( L1195, L1379 ); 
   inv U683 ( L1204, L1380 ); 
   inv U684 ( L1213, L1381 ); 
   inv U685 ( L1222, L1382 ); 
   inv U686 ( L1231, L1383 ); 
   inv U687 ( L1168, L1393 ); 
   inv U688 ( L1177, L1394 ); 
   inv U689 ( L1186, L1395 ); 
   inv U690 ( L1195, L1396 ); 
   inv U691 ( L1204, L1397 ); 
   inv U692 ( L1213, L1398 ); 
   inv U693 ( L1222, L1399 ); 
   inv U694 ( L1231, L1400 ); 
   inv U695 ( L1168, L1410 ); 
   inv U696 ( L1177, L1411 ); 
   inv U697 ( L1186, L1412 ); 
   inv U698 ( L1195, L1413 ); 
   inv U699 ( L1204, L1414 ); 
   inv U700 ( L1213, L1415 ); 
   inv U701 ( L1222, L1416 ); 
   inv U702 ( L1231, L1417 ); 
   inv U703 ( L1168, L1427 ); 
   inv U704 ( L1177, L1428 ); 
   inv U705 ( L1186, L1429 ); 
   inv U706 ( L1195, L1430 ); 
   inv U707 ( L1204, L1431 ); 
   inv U708 ( L1213, L1432 ); 
   inv U709 ( L1222, L1433 ); 
   inv U710 ( L1231, L1434 ); 
   inv U711 ( L1168, L1444 ); 
   inv U712 ( L1177, L1445 ); 
   inv U713 ( L1186, L1446 ); 
   inv U714 ( L1195, L1447 ); 
   inv U715 ( L1204, L1448 ); 
   inv U716 ( L1213, L1449 ); 
   inv U717 ( L1222, L1450 ); 
   inv U718 ( L1231, L1451 ); 
   inv U719 ( L1168, L1461 ); 
   inv U720 ( L1177, L1462 ); 
   inv U721 ( L1186, L1463 ); 
   inv U722 ( L1195, L1464 ); 
   inv U723 ( L1204, L1465 ); 
   inv U724 ( L1213, L1466 ); 
   inv U725 ( L1222, L1467 ); 
   inv U726 ( L1231, L1468 ); 
   inv U727 ( L1168, L1478 ); 
   inv U728 ( L1177, L1479 ); 
   inv U729 ( L1186, L1480 ); 
   inv U730 ( L1195, L1481 ); 
   inv U731 ( L1204, L1482 ); 
   inv U732 ( L1213, L1483 ); 
   inv U733 ( L1222, L1484 ); 
   inv U734 ( L1231, L1485 ); 
   inv U735 ( L1168, L1495 ); 
   inv U736 ( L1177, L1496 ); 
   inv U737 ( L1186, L1497 ); 
   inv U738 ( L1195, L1498 ); 
   inv U739 ( L1204, L1499 ); 
   inv U740 ( L1213, L1500 ); 
   inv U741 ( L1222, L1501 ); 
   inv U742 ( L1231, L1502 ); 
   buffer U743 ( L1874, L1877 ); 
   inv U744 ( L1874, L1880 ); 
   inv U745 ( L1866, L1891 ); 
   and2 U746 ( L986, L1901, L1903 ); 
   buffer U747 ( L1924, L1927 ); 
   inv U748 ( L1924, L1930 ); 
   buffer U749 ( L1975, L1978 ); 
   inv U750 ( L1975, L1981 ); 
   inv U751 ( L1967, L1992 ); 
   buffer U752 ( L2025, L2028 ); 
   inv U753 ( L2025, L2031 ); 
   inv U754 ( L2017, L2042 ); 
   buffer U755 ( L2080, L2085 ); 
   inv U756 ( L2080, L2088 ); 
   inv U757 ( L2072, L2099 ); 
   and2 U758 ( L1014, L2109, L2111 ); 
   buffer U759 ( L2132, L2137 ); 
   inv U760 ( L2132, L2140 ); 
   buffer U761 ( L2185, L2190 ); 
   inv U762 ( L2185, L2193 ); 
   inv U763 ( L2177, L2204 ); 
   buffer U764 ( L2237, L2242 ); 
   inv U765 ( L2237, L2245 ); 
   inv U766 ( L2229, L2256 ); 
   and2 U767 ( L2285, L1862, L2320 ); 
   and2 U768 ( L2289, L1963, L2341 ); 
   and2 U769 ( L2289, L2013, L2354 ); 
   and2 U770 ( L2289, L2068, L2367 ); 
   and2 U771 ( L2298, L2173, L2383 ); 
   and2 U772 ( L2298, L2225, L2391 ); 
   inv U773 ( L2080, L2474 ); 
   inv U774 ( L2132, L2475 ); 
   inv U775 ( L2185, L2476 ); 
   inv U776 ( L2237, L2477 ); 
   and5 U777 ( L2080, L2132, L2185, L2237, L2481, L2482 ); 
   nand2 U778 ( L359, L360, L361 ); 
   inv U779 ( L567, L568 ); 
   or3 U780 ( L614, L616, L617, L618 ); 
   and2 U781 ( L124, L1240, L1248 ); 
   and2 U782 ( L159, L1241, L1249 ); 
   and2 U783 ( L150, L1242, L1250 ); 
   and2 U784 ( L143, L1243, L1251 ); 
   and2 U785 ( L137, L1244, L1252 ); 
   and2 U786 ( L132, L1245, L1253 ); 
   and2 U787 ( L128, L1246, L1254 ); 
   and2 U788 ( L125, L1247, L1255 ); 
   and2 U789 ( L125, L1257, L1265 ); 
   and2 U790 ( L432, L1258, L1266 ); 
   and2 U791 ( L159, L1259, L1267 ); 
   and2 U792 ( L150, L1260, L1268 ); 
   and2 U793 ( L143, L1261, L1269 ); 
   and2 U794 ( L137, L1262, L1270 ); 
   and2 U795 ( L132, L1263, L1271 ); 
   and2 U796 ( L128, L1264, L1272 ); 
   and2 U797 ( L128, L1274, L1282 ); 
   and2 U798 ( L447, L1275, L1283 ); 
   and2 U799 ( L432, L1276, L1284 ); 
   and2 U800 ( L159, L1277, L1285 ); 
   and2 U801 ( L150, L1278, L1286 ); 
   and2 U802 ( L143, L1279, L1287 ); 
   and2 U803 ( L137, L1280, L1288 ); 
   and2 U804 ( L132, L1281, L1289 ); 
   and2 U805 ( L132, L1291, L1299 ); 
   and2 U806 ( L467, L1292, L1300 ); 
   and2 U807 ( L447, L1293, L1301 ); 
   and2 U808 ( L432, L1294, L1302 ); 
   and2 U809 ( L159, L1295, L1303 ); 
   and2 U810 ( L150, L1296, L1304 ); 
   and2 U811 ( L143, L1297, L1305 ); 
   and2 U812 ( L137, L1298, L1306 ); 
   and2 U813 ( L137, L1308, L1316 ); 
   and2 U814 ( L483, L1309, L1317 ); 
   and2 U815 ( L467, L1310, L1318 ); 
   and2 U816 ( L447, L1311, L1319 ); 
   and2 U817 ( L432, L1312, L1320 ); 
   and2 U818 ( L159, L1313, L1321 ); 
   and2 U819 ( L150, L1314, L1322 ); 
   and2 U820 ( L143, L1315, L1323 ); 
   and2 U821 ( L143, L1325, L1333 ); 
   and2 U822 ( L492, L1326, L1334 ); 
   and2 U823 ( L483, L1327, L1335 ); 
   and2 U824 ( L467, L1328, L1336 ); 
   and2 U825 ( L447, L1329, L1337 ); 
   and2 U826 ( L432, L1330, L1338 ); 
   and2 U827 ( L159, L1331, L1339 ); 
   and2 U828 ( L150, L1332, L1340 ); 
   and2 U829 ( L150, L1342, L1350 ); 
   and2 U830 ( L504, L1343, L1351 ); 
   and2 U831 ( L492, L1344, L1352 ); 
   and2 U832 ( L483, L1345, L1353 ); 
   and2 U833 ( L467, L1346, L1354 ); 
   and2 U834 ( L447, L1347, L1355 ); 
   and2 U835 ( L432, L1348, L1356 ); 
   and2 U836 ( L159, L1349, L1357 ); 
   and2 U837 ( L159, L1359, L1367 ); 
   and2 U838 ( L517, L1360, L1368 ); 
   and2 U839 ( L504, L1361, L1369 ); 
   and2 U840 ( L492, L1362, L1370 ); 
   and2 U841 ( L483, L1363, L1371 ); 
   and2 U842 ( L467, L1364, L1372 ); 
   and2 U843 ( L447, L1365, L1373 ); 
   and2 U844 ( L432, L1366, L1374 ); 
   and2 U845 ( L283, L1376, L1384 ); 
   and2 U846 ( L447, L1377, L1385 ); 
   and2 U847 ( L467, L1378, L1386 ); 
   and2 U848 ( L483, L1379, L1387 ); 
   and2 U849 ( L492, L1380, L1388 ); 
   and2 U850 ( L504, L1381, L1389 ); 
   and2 U851 ( L517, L1382, L1390 ); 
   and2 U852 ( L530, L1383, L1391 ); 
   and2 U853 ( L294, L1393, L1401 ); 
   and2 U854 ( L467, L1394, L1402 ); 
   and2 U855 ( L483, L1395, L1403 ); 
   and2 U856 ( L492, L1396, L1404 ); 
   and2 U857 ( L504, L1397, L1405 ); 
   and2 U858 ( L517, L1398, L1406 ); 
   and2 U859 ( L530, L1399, L1407 ); 
   and2 U860 ( L283, L1400, L1408 ); 
   and2 U861 ( L303, L1410, L1418 ); 
   and2 U862 ( L483, L1411, L1419 ); 
   and2 U863 ( L492, L1412, L1420 ); 
   and2 U864 ( L504, L1413, L1421 ); 
   and2 U865 ( L517, L1414, L1422 ); 
   and2 U866 ( L530, L1415, L1423 ); 
   and2 U867 ( L283, L1416, L1424 ); 
   and2 U868 ( L294, L1417, L1425 ); 
   and2 U869 ( L311, L1427, L1435 ); 
   and2 U870 ( L492, L1428, L1436 ); 
   and2 U871 ( L504, L1429, L1437 ); 
   and2 U872 ( L517, L1430, L1438 ); 
   and2 U873 ( L530, L1431, L1439 ); 
   and2 U874 ( L283, L1432, L1440 ); 
   and2 U875 ( L294, L1433, L1441 ); 
   and2 U876 ( L303, L1434, L1442 ); 
   and2 U877 ( L317, L1444, L1452 ); 
   and2 U878 ( L504, L1445, L1453 ); 
   and2 U879 ( L517, L1446, L1454 ); 
   and2 U880 ( L530, L1447, L1455 ); 
   and2 U881 ( L283, L1448, L1456 ); 
   and2 U882 ( L294, L1449, L1457 ); 
   and2 U883 ( L303, L1450, L1458 ); 
   and2 U884 ( L311, L1451, L1459 ); 
   and2 U885 ( L322, L1461, L1469 ); 
   and2 U886 ( L517, L1462, L1470 ); 
   and2 U887 ( L530, L1463, L1471 ); 
   and2 U888 ( L283, L1464, L1472 ); 
   and2 U889 ( L294, L1465, L1473 ); 
   and2 U890 ( L303, L1466, L1474 ); 
   and2 U891 ( L311, L1467, L1475 ); 
   and2 U892 ( L317, L1468, L1476 ); 
   and2 U893 ( L326, L1478, L1486 ); 
   and2 U894 ( L530, L1479, L1487 ); 
   and2 U895 ( L283, L1480, L1488 ); 
   and2 U896 ( L294, L1481, L1489 ); 
   and2 U897 ( L303, L1482, L1490 ); 
   and2 U898 ( L311, L1483, L1491 ); 
   and2 U899 ( L317, L1484, L1492 ); 
   and2 U900 ( L322, L1485, L1493 ); 
   and2 U901 ( L329, L1495, L1503 ); 
   and2 U902 ( L283, L1496, L1504 ); 
   and2 U903 ( L294, L1497, L1505 ); 
   and2 U904 ( L303, L1498, L1506 ); 
   and2 U905 ( L311, L1499, L1507 ); 
   and2 U906 ( L317, L1500, L1508 ); 
   and2 U907 ( L322, L1501, L1509 ); 
   and2 U908 ( L326, L1502, L1510 ); 
   and5 U909 ( L2474, L2475, L2476, L2477, L2478, L2483 ); 
   buffer U910 ( L597, L600 ); 
   and2 U911 ( L568, L660, L661 ); 
   and2 U912 ( L597, L665, L669 ); 
   and2 U913 ( L591, L678, L679 ); 
   nor8 U914 ( L1248, L1249, L1250, L1251, L1252, L1253, L1254, L1255, L1256 ); 
   nor8 U915 ( L1265, L1266, L1267, L1268, L1269, L1270, L1271, L1272, L1273 ); 
   nor8 U916 ( L1282, L1283, L1284, L1285, L1286, L1287, L1288, L1289, L1290 ); 
   nor8 U917 ( L1299, L1300, L1301, L1302, L1303, L1304, L1305, L1306, L1307 ); 
   nor8 U918 ( L1316, L1317, L1318, L1319, L1320, L1321, L1322, L1323, L1324 ); 
   nor8 U919 ( L1333, L1334, L1335, L1336, L1337, L1338, L1339, L1340, L1341 ); 
   nor8 U920 ( L1350, L1351, L1352, L1353, L1354, L1355, L1356, L1357, L1358 ); 
   nor8 U921 ( L1367, L1368, L1369, L1370, L1371, L1372, L1373, L1374, L1375 ); 
   nor8 U922 ( L1384, L1385, L1386, L1387, L1388, L1389, L1390, L1391, L1392 ); 
   nor8 U923 ( L1401, L1402, L1403, L1404, L1405, L1406, L1407, L1408, L1409 ); 
   nor8 U924 ( L1418, L1419, L1420, L1421, L1422, L1423, L1424, L1425, L1426 ); 
   nor8 U925 ( L1435, L1436, L1437, L1438, L1439, L1440, L1441, L1442, L1443 ); 
   nor8 U926 ( L1452, L1453, L1454, L1455, L1456, L1457, L1458, L1459, L1460 ); 
   nor8 U927 ( L1469, L1470, L1471, L1472, L1473, L1474, L1475, L1476, L1477 ); 
   nor8 U928 ( L1486, L1487, L1488, L1489, L1490, L1491, L1492, L1493, L1494 ); 
   nor8 U929 ( L1503, L1504, L1505, L1506, L1507, L1508, L1509, L1510, L1511 ); 
   and2 U930 ( L618, L1647, L1652 ); 
   and3 U931 ( L169, L1862, L1877, L1883 ); 
   and3 U932 ( L179, L1862, L1880, L1886 ); 
   and3 U933 ( L190, L1866, L1880, L1889 ); 
   and3 U934 ( L200, L1866, L1877, L1890 ); 
   or3 U935 ( L1903, L1906, L1909, L1912 ); 
   nor3 U936 ( L1903, L1906, L1909, L1916 ); 
   and3 U937 ( L169, L1963, L1978, L1984 ); 
   and3 U938 ( L179, L1963, L1981, L1987 ); 
   and3 U939 ( L190, L1967, L1981, L1990 ); 
   and3 U940 ( L200, L1967, L1978, L1991 ); 
   and3 U941 ( L169, L2013, L2028, L2034 ); 
   and3 U942 ( L179, L2013, L2031, L2037 ); 
   and3 U943 ( L190, L2017, L2031, L2040 ); 
   and3 U944 ( L200, L2017, L2028, L2041 ); 
   and3 U945 ( L169, L2068, L2085, L2091 ); 
   and3 U946 ( L179, L2068, L2088, L2094 ); 
   and3 U947 ( L190, L2072, L2088, L2097 ); 
   and3 U948 ( L200, L2072, L2085, L2098 ); 
   or3 U949 ( L2111, L2114, L2117, L2120 ); 
   nor3 U950 ( L2111, L2114, L2117, L2124 ); 
   and3 U951 ( L169, L2173, L2190, L2196 ); 
   and3 U952 ( L179, L2173, L2193, L2199 ); 
   and3 U953 ( L190, L2177, L2193, L2202 ); 
   and3 U954 ( L200, L2177, L2190, L2203 ); 
   and3 U955 ( L169, L2225, L2242, L2248 ); 
   and3 U956 ( L179, L2225, L2245, L2251 ); 
   and3 U957 ( L190, L2229, L2245, L2254 ); 
   and3 U958 ( L200, L2229, L2242, L2255 ); 
   or2 U959 ( L2482, L2483, L2484 ); 
   buffer U960 ( L571, L2991 ); 
   buffer U961 ( L579, L2994 ); 
   buffer U962 ( L571, L2999 ); 
   buffer U963 ( L579, L3002 ); 
   buffer U964 ( L591, L3063 ); 
   buffer U965 ( L591, L3071 ); 
   buffer U966 ( L2320, L3124 ); 
   buffer U967 ( L2320, L3134 ); 
   buffer U968 ( L2341, L3158 ); 
   buffer U969 ( L2341, L3166 ); 
   buffer U970 ( L2354, L3174 ); 
   buffer U971 ( L2354, L3182 ); 
   buffer U972 ( L2367, L3190 ); 
   buffer U973 ( L2367, L3200 ); 
   buffer U974 ( L2383, L3224 ); 
   buffer U975 ( L2383, L3232 ); 
   buffer U976 ( L2391, L3240 ); 
   buffer U977 ( L2391, L3248 ); 
   nor2 U978 ( L661, L662, L663 ); 
   or3 U979 ( L669, L671, L672, L673 ); 
   nor2 U980 ( L679, L680, L681 ); 
   and2 U981 ( L1256, L1533, L1536 ); 
   and2 U982 ( L1392, L1534, L1537 ); 
   and2 U983 ( L1273, L1581, L1582 ); 
   and2 U984 ( L1409, L1512, L1583 ); 
   and2 U985 ( L1290, L1585, L1586 ); 
   and2 U986 ( L1426, L1512, L1587 ); 
   and2 U987 ( L1307, L1589, L1590 ); 
   and2 U988 ( L1443, L1512, L1591 ); 
   and2 U989 ( L1324, L1593, L1594 ); 
   and2 U990 ( L1460, L1512, L1595 ); 
   and2 U991 ( L1341, L1597, L1598 ); 
   and2 U992 ( L1477, L1512, L1599 ); 
   and2 U993 ( L1358, L1601, L1602 ); 
   and2 U994 ( L1494, L1512, L1603 ); 
   and2 U995 ( L1375, L1605, L1606 ); 
   and2 U996 ( L1511, L1512, L1607 ); 
   or3 U997 ( L1889, L1890, L1891, L1894 ); 
   or3 U998 ( L1990, L1991, L1992, L1997 ); 
   or3 U999 ( L2040, L2041, L2042, L2047 ); 
   or3 U1000 ( L2097, L2098, L2099, L2102 ); 
   or3 U1001 ( L2202, L2203, L2204, L2209 ); 
   or3 U1002 ( L2254, L2255, L2256, L2261 ); 
   and2 U1003 ( L2484, L2488, L2489 ); 
   inv U1004 ( L2999, L3005 ); 
   inv U1005 ( L3002, L3006 ); 
   inv U1006 ( L3071, L3077 ); 
   inv U1007 ( L3063, L3069 ); 
   inv U1008 ( L2991, L2997 ); 
   inv U1009 ( L2994, L2998 ); 
   and2 U1010 ( L681, L683, L689 ); 
   and2 U1011 ( L663, L694, L700 ); 
   or3 U1012 ( L1536, L1537, L1538, L1539 ); 
   or2 U1013 ( L1582, L1583, L1584 ); 
   or2 U1014 ( L1586, L1587, L1588 ); 
   or2 U1015 ( L1590, L1591, L1592 ); 
   or2 U1016 ( L1594, L1595, L1596 ); 
   or2 U1017 ( L1598, L1599, L1600 ); 
   or2 U1018 ( L1602, L1603, L1604 ); 
   or2 U1019 ( L1606, L1607, L1608 ); 
   and2 U1020 ( L673, L1656, L1661 ); 
   or2 U1021 ( L1883, L1886, L1892 ); 
   nor2 U1022 ( L1883, L1886, L1893 ); 
   and3 U1023 ( L169, L1912, L1927, L1933 ); 
   and3 U1024 ( L179, L1912, L1930, L1936 ); 
   and3 U1025 ( L190, L1916, L1930, L1939 ); 
   and3 U1026 ( L200, L1916, L1927, L1940 ); 
   inv U1027 ( L1916, L1941 ); 
   or2 U1028 ( L1984, L1987, L1993 ); 
   nor2 U1029 ( L1984, L1987, L1996 ); 
   or2 U1030 ( L2034, L2037, L2043 ); 
   nor2 U1031 ( L2034, L2037, L2046 ); 
   or2 U1032 ( L2091, L2094, L2100 ); 
   nor2 U1033 ( L2091, L2094, L2101 ); 
   and3 U1034 ( L169, L2120, L2137, L2143 ); 
   and3 U1035 ( L179, L2120, L2140, L2146 ); 
   and3 U1036 ( L190, L2124, L2140, L2149 ); 
   and3 U1037 ( L200, L2124, L2137, L2150 ); 
   inv U1038 ( L2124, L2151 ); 
   or2 U1039 ( L2196, L2199, L2205 ); 
   nor2 U1040 ( L2196, L2199, L2208 ); 
   or2 U1041 ( L2248, L2251, L2257 ); 
   nor2 U1042 ( L2248, L2251, L2260 ); 
   inv U1043 ( L3134, L3138 ); 
   and2 U1044 ( L2285, L1912, L2328 ); 
   inv U1045 ( L3158, L3162 ); 
   inv U1046 ( L3166, L3170 ); 
   inv U1047 ( L3174, L3178 ); 
   inv U1048 ( L3182, L3186 ); 
   inv U1049 ( L3200, L3204 ); 
   and2 U1050 ( L2298, L2120, L2375 ); 
   inv U1051 ( L3232, L3236 ); 
   inv U1052 ( L3240, L3244 ); 
   inv U1053 ( L3248, L3252 ); 
   inv U1054 ( L3224, L3228 ); 
   buffer U1055 ( L600, L3066 ); 
   buffer U1056 ( L600, L3074 ); 
   inv U1057 ( L3124, L3128 ); 
   inv U1058 ( L3190, L3194 ); 
   nand2 U1059 ( L2994, L2997, L619 ); 
   nand2 U1060 ( L2991, L2998, L620 ); 
   nand2 U1061 ( L3002, L3005, L582 ); 
   nand2 U1062 ( L2999, L3006, L583 ); 
   or3 U1063 ( L689, L690, L691, L692 ); 
   or3 U1064 ( L700, L701, L702, L703 ); 
   and2 U1065 ( L1539, L1609, L1612 ); 
   and2 U1066 ( L1584, L1618, L1621 ); 
   and2 U1067 ( L1588, L1627, L1630 ); 
   and2 U1068 ( L1592, L1636, L1639 ); 
   and2 U1069 ( L1596, L1645, L1648 ); 
   and2 U1070 ( L1600, L1654, L1657 ); 
   and2 U1071 ( L1604, L1663, L1666 ); 
   and2 U1072 ( L1608, L1672, L1675 ); 
   and2 U1073 ( L1893, L1894, L1895 ); 
   or3 U1074 ( L1939, L1940, L1941, L1946 ); 
   and2 U1075 ( L1996, L1997, L1998 ); 
   and2 U1076 ( L2046, L2047, L2048 ); 
   and2 U1077 ( L2101, L2102, L2103 ); 
   or3 U1078 ( L2149, L2150, L2151, L2156 ); 
   and2 U1079 ( L2208, L2209, L2210 ); 
   and2 U1080 ( L2260, L2261, L2262 ); 
   inv U1081 ( L1892, L2271 ); 
   inv U1082 ( L2100, L2311 ); 
   nand2 U1083 ( L619, L620, L356 ); 
   nand2 U1084 ( L582, L583, L357 ); 
   nand2 U1085 ( L3074, L3077, L603 ); 
   inv U1086 ( L3074, L3078 ); 
   nand2 U1087 ( L3066, L3069, L606 ); 
   inv U1088 ( L3066, L3070 ); 
   and2 U1089 ( L703, L1665, L1670 ); 
   and2 U1090 ( L692, L1674, L1679 ); 
   or2 U1091 ( L1933, L1936, L1942 ); 
   nor2 U1092 ( L1933, L1936, L1945 ); 
   or2 U1093 ( L2143, L2146, L2152 ); 
   nor2 U1094 ( L2143, L2146, L2155 ); 
   and2 U1095 ( L1993, L2293, L2445 ); 
   and2 U1096 ( L2043, L2293, L2448 ); 
   and2 U1097 ( L2205, L2302, L2455 ); 
   and2 U1098 ( L2257, L2302, L2458 ); 
   buffer U1099 ( L2328, L3142 ); 
   buffer U1100 ( L2328, L3150 ); 
   buffer U1101 ( L2375, L3208 ); 
   buffer U1102 ( L2375, L3216 ); 
   nand2 U1103 ( L356, L357, L358 ); 
   nand2 U1104 ( L3071, L3078, L604 ); 
   nand2 U1105 ( L3063, L3070, L607 ); 
   and2 U1106 ( L1945, L1946, L1947 ); 
   and2 U1107 ( L2155, L2156, L2157 ); 
   buffer U1108 ( L1895, L2317 ); 
   buffer U1109 ( L1998, L2338 ); 
   buffer U1110 ( L2048, L2351 ); 
   buffer U1111 ( L2103, L2364 ); 
   buffer U1112 ( L2210, L2380 ); 
   buffer U1113 ( L2262, L2388 ); 
   nand2 U1114 ( L603, L604, L605 ); 
   nand2 U1115 ( L606, L607, L608 ); 
   nand2 U1116 ( L1895, L1942, L2272 ); 
   nand2 U1117 ( L2103, L2152, L2312 ); 
   inv U1118 ( L3142, L3146 ); 
   inv U1119 ( L3150, L3154 ); 
   inv U1120 ( L3216, L3220 ); 
   inv U1121 ( L3208, L3212 ); 
   and2 U1122 ( L1942, L2288, L2444 ); 
   buffer U1123 ( L2448, L2451 ); 
   and2 U1124 ( L2152, L2293, L2454 ); 
   buffer U1125 ( L2458, L2461 ); 
   inv U1126 ( L2445, L2530 ); 
   buffer U1127 ( L2458, L3323 ); 
   inv U1128 ( L605, L349 ); 
   inv U1129 ( L608, L350 ); 
   and4 U1130 ( L1895, L1947, L1998, L2048, L2265 ); 
   nand3 U1131 ( L1895, L1947, L1993, L2273 ); 
   nand4 U1132 ( L2043, L1947, L1998, L1895, L2274 ); 
   and4 U1133 ( L2103, L2157, L2210, L2262, L2309 ); 
   nand3 U1134 ( L2103, L2157, L2205, L2313 ); 
   nand4 U1135 ( L2257, L2157, L2210, L2103, L2314 ); 
   buffer U1136 ( L1947, L2325 ); 
   buffer U1137 ( L2157, L2372 ); 
   inv U1138 ( L2444, L2523 ); 
   inv U1139 ( L2454, L2533 ); 
   buffer U1140 ( L2317, L3121 ); 
   buffer U1141 ( L2317, L3131 ); 
   buffer U1142 ( L2338, L3155 ); 
   buffer U1143 ( L2338, L3163 ); 
   buffer U1144 ( L2351, L3171 ); 
   buffer U1145 ( L2351, L3179 ); 
   buffer U1146 ( L2364, L3187 ); 
   buffer U1147 ( L2364, L3197 ); 
   buffer U1148 ( L2380, L3221 ); 
   buffer U1149 ( L2380, L3229 ); 
   buffer U1150 ( L2388, L3237 ); 
   buffer U1151 ( L2388, L3245 ); 
   nand2 U1152 ( L349, L350, L351 ); 
   nand4 U1153 ( L2271, L2272, L2273, L2274, L2275 ); 
   nand4 U1154 ( L2311, L2312, L2313, L2314, L2315 ); 
   inv U1155 ( L3323, L3329 ); 
   and2 U1156 ( L2309, L2265, L372 ); 
   nand2 U1157 ( L3131, L3138, L2324 ); 
   nand2 U1158 ( L3163, L3170, L2350 ); 
   nand2 U1159 ( L3179, L3186, L2363 ); 
   nand2 U1160 ( L3197, L3204, L2371 ); 
   nand2 U1161 ( L3229, L3236, L2387 ); 
   nand2 U1162 ( L3245, L3252, L2400 ); 
   buffer U1163 ( L2265, L2268 ); 
   inv U1164 ( L3131, L3137 ); 
   inv U1165 ( L3155, L3161 ); 
   nand2 U1166 ( L3155, L3162, L2345 ); 
   inv U1167 ( L3163, L3169 ); 
   inv U1168 ( L3171, L3177 ); 
   nand2 U1169 ( L3171, L3178, L2358 ); 
   inv U1170 ( L3179, L3185 ); 
   inv U1171 ( L3197, L3203 ); 
   inv U1172 ( L3229, L3235 ); 
   inv U1173 ( L3237, L3243 ); 
   nand2 U1174 ( L3237, L3244, L2395 ); 
   inv U1175 ( L3245, L3251 ); 
   inv U1176 ( L3221, L3227 ); 
   nand2 U1177 ( L3221, L3228, L2432 ); 
   and2 U1178 ( L2309, L2485, L2490 ); 
   inv U1179 ( L3121, L3127 ); 
   nand2 U1180 ( L3121, L3128, L3130 ); 
   buffer U1181 ( L2325, L3139 ); 
   buffer U1182 ( L2325, L3147 ); 
   inv U1183 ( L3187, L3193 ); 
   nand2 U1184 ( L3187, L3194, L3196 ); 
   buffer U1185 ( L2372, L3205 ); 
   buffer U1186 ( L2372, L3213 ); 
   nand2 U1187 ( L2265, L2315, L2307 ); 
   inv U1188 ( L2275, L2308 ); 
   nand2 U1189 ( L3134, L3137, L2323 ); 
   nand2 U1190 ( L3166, L3169, L2349 ); 
   nand2 U1191 ( L3182, L3185, L2362 ); 
   nand2 U1192 ( L3200, L3203, L2370 ); 
   nand2 U1193 ( L3232, L3235, L2386 ); 
   nand2 U1194 ( L3248, L3251, L2399 ); 
   nand2 U1195 ( L3158, L3161, L2344 ); 
   nand2 U1196 ( L3174, L3177, L2357 ); 
   nand2 U1197 ( L3240, L3243, L2394 ); 
   nand2 U1198 ( L3224, L3227, L2431 ); 
   and2 U1199 ( L2315, L2302, L2464 ); 
   or2 U1200 ( L2489, L2490, L2491 ); 
   nand2 U1201 ( L3124, L3127, L3129 ); 
   nand2 U1202 ( L3190, L3193, L3195 ); 
   and2 U1203 ( L2307, L2308, L368 ); 
   nand2 U1204 ( L2323, L2324, L1615 ); 
   nand2 U1205 ( L3147, L3154, L2337 ); 
   nand2 U1206 ( L2349, L2350, L1633 ); 
   nand2 U1207 ( L2362, L2363, L1642 ); 
   nand2 U1208 ( L2370, L2371, L1651 ); 
   nand2 U1209 ( L3213, L3220, L2379 ); 
   nand2 U1210 ( L2386, L2387, L1669 ); 
   nand2 U1211 ( L2399, L2400, L1678 ); 
   inv U1212 ( L3139, L3145 ); 
   nand2 U1213 ( L3139, L3146, L2332 ); 
   inv U1214 ( L3147, L3153 ); 
   nand2 U1215 ( L2344, L2345, L2346 ); 
   nand2 U1216 ( L2357, L2358, L2359 ); 
   inv U1217 ( L3213, L3219 ); 
   nand2 U1218 ( L2394, L2395, L2396 ); 
   inv U1219 ( L3205, L3211 ); 
   nand2 U1220 ( L3205, L3212, L2425 ); 
   nand2 U1221 ( L2431, L2432, L2433 ); 
   nand2 U1222 ( L3129, L3130, L3272 ); 
   nand2 U1223 ( L3195, L3196, L3308 ); 
   inv U1224 ( L368, L369 ); 
   inv U1225 ( L1615, L1613 ); 
   nand2 U1226 ( L3150, L3153, L2336 ); 
   inv U1227 ( L1633, L1631 ); 
   inv U1228 ( L1642, L1640 ); 
   inv U1229 ( L1651, L1649 ); 
   nand2 U1230 ( L3216, L3219, L2378 ); 
   inv U1231 ( L1669, L1667 ); 
   inv U1232 ( L1678, L1676 ); 
   nand2 U1233 ( L3142, L3145, L2331 ); 
   nand2 U1234 ( L3208, L3211, L2424 ); 
   buffer U1235 ( L2464, L2467 ); 
   buffer U1236 ( L2491, L2495 ); 
   buffer U1237 ( L2464, L3295 ); 
   and2 U1238 ( L330, L2491, L3374 ); 
   and2 U1239 ( L1613, L1610, L1614 ); 
   nand2 U1240 ( L2336, L2337, L1624 ); 
   and2 U1241 ( L1631, L1628, L1632 ); 
   and2 U1242 ( L1640, L1637, L1641 ); 
   and2 U1243 ( L1649, L1646, L1650 ); 
   nand2 U1244 ( L2378, L2379, L1660 ); 
   and2 U1245 ( L1667, L1664, L1668 ); 
   and2 U1246 ( L1676, L1673, L1677 ); 
   nand2 U1247 ( L2331, L2332, L2333 ); 
   buffer U1248 ( L2346, L2406 ); 
   buffer U1249 ( L2346, L2409 ); 
   buffer U1250 ( L2359, L2415 ); 
   buffer U1251 ( L2359, L2419 ); 
   nand2 U1252 ( L2424, L2425, L2426 ); 
   buffer U1253 ( L2396, L2439 ); 
   and2 U1254 ( L2433, L2461, L2518 ); 
   inv U1255 ( L3272, L3276 ); 
   inv U1256 ( L3308, L3312 ); 
   and2 U1257 ( L330, L2396, L2612 ); 
   buffer U1258 ( L2433, L3326 ); 
   nor3 U1259 ( L1612, L1614, L1616, L1617 ); 
   inv U1260 ( L1624, L1622 ); 
   nor3 U1261 ( L1630, L1632, L1634, L1635 ); 
   nor3 U1262 ( L1639, L1641, L1643, L1644 ); 
   nor3 U1263 ( L1648, L1650, L1652, L1653 ); 
   inv U1264 ( L1660, L1658 ); 
   nor3 U1265 ( L1666, L1668, L1670, L1671 ); 
   nor3 U1266 ( L1675, L1677, L1679, L1680 ); 
   and2 U1267 ( L2467, L2268, L2500 ); 
   and2 U1268 ( L2495, L2268, L2505 ); 
   or2 U1269 ( L2455, L2518, L2519 ); 
   inv U1270 ( L3374, L3378 ); 
   inv U1271 ( L2467, L2642 ); 
   buffer U1272 ( L2467, L2645 ); 
   inv U1273 ( L3295, L3301 ); 
   and2 U1274 ( L1622, L1619, L1623 ); 
   and2 U1275 ( L1658, L1655, L1659 ); 
   buffer U1276 ( L2333, L2401 ); 
   or2 U1277 ( L2275, L2500, L2501 ); 
   and3 U1278 ( L2495, L2419, L2409, L2511 ); 
   and2 U1279 ( L2495, L2415, L2512 ); 
   and3 U1280 ( L2439, L2433, L2426, L2513 ); 
   and2 U1281 ( L2439, L2433, L2514 ); 
   and2 U1282 ( L2467, L2415, L2517 ); 
   nand2 U1283 ( L2409, L2451, L2531 ); 
   nand3 U1284 ( L2409, L2419, L2467, L2532 ); 
   nand2 U1285 ( L2426, L2455, L2534 ); 
   nand3 U1286 ( L2426, L2433, L2461, L2535 ); 
   nand2 U1287 ( L3326, L3329, L2607 ); 
   inv U1288 ( L3326, L3330 ); 
   and3 U1289 ( L330, L2491, L2642, L2643 ); 
   and2 U1290 ( L1617, L2680, L2687 ); 
   and2 U1291 ( L1635, L2718, L2725 ); 
   and2 U1292 ( L1644, L2735, L2742 ); 
   and2 U1293 ( L1653, L2753, L2760 ); 
   and2 U1294 ( L1671, L2787, L2794 ); 
   and2 U1295 ( L1680, L2804, L2811 ); 
   buffer U1296 ( L2333, L3280 ); 
   buffer U1297 ( L2409, L3290 ); 
   buffer U1298 ( L2415, L3298 ); 
   buffer U1299 ( L2426, L3316 ); 
   buffer U1300 ( L2612, L3406 ); 
   buffer U1301 ( L2612, L3414 ); 
   buffer U1302 ( L2439, L3422 ); 
   nor3 U1303 ( L1621, L1623, L1625, L1626 ); 
   nor3 U1304 ( L1657, L1659, L1661, L1662 ); 
   and2 U1305 ( L330, L2512, L2567 ); 
   and2 U1306 ( L330, L2513, L2589 ); 
   nand2 U1307 ( L3323, L3330, L2608 ); 
   buffer U1308 ( L2519, L2654 ); 
   buffer U1309 ( L2505, L3253 ); 
   nand3 U1310 ( L2530, L2531, L2532, L3277 ); 
   or2 U1311 ( L2448, L2517, L3287 ); 
   nand3 U1312 ( L2533, L2534, L2535, L3305 ); 
   buffer U1313 ( L2519, L3313 ); 
   and2 U1314 ( L330, L2511, L3350 ); 
   or2 U1315 ( L2643, L2645, L932 ); 
   and4 U1316 ( L2495, L2401, L2409, L2419, L2508 ); 
   nand2 U1317 ( L2401, L2445, L2524 ); 
   nand3 U1318 ( L2401, L2406, L2451, L2525 ); 
   nand4 U1319 ( L2401, L2406, L2419, L2467, L2526 ); 
   inv U1320 ( L3290, L3294 ); 
   nand2 U1321 ( L2607, L2608, L2609 ); 
   inv U1322 ( L3406, L3410 ); 
   inv U1323 ( L3414, L3418 ); 
   nand2 U1324 ( L3422, L3425, L2624 ); 
   inv U1325 ( L3422, L3426 ); 
   buffer U1326 ( L2501, L2629 ); 
   nor2 U1327 ( L2643, L2645, L2647 ); 
   and2 U1328 ( L1626, L2699, L2706 ); 
   and2 U1329 ( L1662, L2770, L2777 ); 
   buffer U1330 ( L2501, L3264 ); 
   inv U1331 ( L3280, L3284 ); 
   inv U1332 ( L3298, L3302 ); 
   nand2 U1333 ( L3298, L3301, L3303 ); 
   inv U1334 ( L3316, L3320 ); 
   and2 U1335 ( L330, L2514, L3398 ); 
   inv U1336 ( L2654, L2657 ); 
   and2 U1337 ( L2519, L2654, L398 ); 
   and2 U1338 ( L932, L927, L933 ); 
   nand4 U1339 ( L2523, L2524, L2525, L2526, L2527 ); 
   inv U1340 ( L3253, L3259 ); 
   inv U1341 ( L3350, L3354 ); 
   inv U1342 ( L3287, L3293 ); 
   nand2 U1343 ( L3287, L3294, L2563 ); 
   inv U1344 ( L3305, L3311 ); 
   nand2 U1345 ( L3305, L3312, L2585 ); 
   nand2 U1346 ( L3419, L3426, L2625 ); 
   inv U1347 ( L3277, L3283 ); 
   nand2 U1348 ( L3277, L3284, L3286 ); 
   nand2 U1349 ( L3295, L3302, L3304 ); 
   inv U1350 ( L3313, L3319 ); 
   nand2 U1351 ( L3313, L3320, L3322 ); 
   buffer U1352 ( L2567, L3358 ); 
   buffer U1353 ( L2567, L3366 ); 
   buffer U1354 ( L2589, L3382 ); 
   buffer U1355 ( L2589, L3390 ); 
   and3 U1356 ( L330, L2514, L2657, L397 ); 
   and2 U1357 ( L330, L2508, L2544 ); 
   nand2 U1358 ( L3290, L3293, L2562 ); 
   nand2 U1359 ( L3308, L3311, L2584 ); 
   inv U1360 ( L3398, L3402 ); 
   nand2 U1361 ( L2624, L2625, L2626 ); 
   inv U1362 ( L2629, L2632 ); 
   and2 U1363 ( L2501, L2629, L2634 ); 
   buffer U1364 ( L2647, L2650 ); 
   inv U1365 ( L3264, L3268 ); 
   buffer U1366 ( L2508, L3256 ); 
   nand2 U1367 ( L3280, L3283, L3285 ); 
   nand2 U1368 ( L3316, L3319, L3321 ); 
   nand2 U1369 ( L3303, L3304, L3371 ); 
   buffer U1370 ( L2609, L3403 ); 
   buffer U1371 ( L2609, L3411 ); 
   or3 U1372 ( L929, L933, L938, L362 ); 
   nor3 U1373 ( L929, L933, L938, L1030 ); 
   or2 U1374 ( L397, L398, L399 ); 
   nand2 U1375 ( L2562, L2563, L2564 ); 
   inv U1376 ( L3358, L3362 ); 
   inv U1377 ( L3366, L3370 ); 
   nand2 U1378 ( L2584, L2585, L2586 ); 
   inv U1379 ( L3382, L3386 ); 
   inv U1380 ( L3390, L3394 ); 
   and3 U1381 ( L330, L2505, L2632, L2633 ); 
   buffer U1382 ( L2527, L3261 ); 
   buffer U1383 ( L2527, L3269 ); 
   nand2 U1384 ( L3285, L3286, L3347 ); 
   nand2 U1385 ( L3321, L3322, L3395 ); 
   inv U1386 ( L1030, L363 ); 
   nand2 U1387 ( L3256, L3259, L2536 ); 
   inv U1388 ( L3256, L3260 ); 
   inv U1389 ( L3371, L3377 ); 
   nand2 U1390 ( L3371, L3378, L2580 ); 
   inv U1391 ( L3403, L3409 ); 
   nand2 U1392 ( L3403, L3410, L2616 ); 
   inv U1393 ( L3411, L3417 ); 
   nand2 U1394 ( L3411, L3418, L2622 ); 
   nor2 U1395 ( L2633, L2634, L2635 ); 
   and2 U1396 ( L2626, L2802, L2805 ); 
   and2 U1397 ( L2626, L2803, L2808 ); 
   buffer U1398 ( L2544, L3334 ); 
   buffer U1399 ( L2544, L3342 ); 
   buffer U1400 ( L2650, L3454 ); 
   and2 U1401 ( L362, L363, L364 ); 
   nand2 U1402 ( L3253, L3260, L2537 ); 
   inv U1403 ( L3269, L3275 ); 
   nand2 U1404 ( L3269, L3276, L2540 ); 
   inv U1405 ( L3347, L3353 ); 
   nand2 U1406 ( L3347, L3354, L2557 ); 
   nand2 U1407 ( L3374, L3377, L2579 ); 
   inv U1408 ( L3395, L3401 ); 
   nand2 U1409 ( L3395, L3402, L2602 ); 
   nand2 U1410 ( L3406, L3409, L2615 ); 
   nand2 U1411 ( L3414, L3417, L2621 ); 
   inv U1412 ( L3261, L3267 ); 
   nand2 U1413 ( L3261, L3268, L3112 ); 
   buffer U1414 ( L2564, L3355 ); 
   buffer U1415 ( L2564, L3363 ); 
   buffer U1416 ( L2586, L3379 ); 
   buffer U1417 ( L2586, L3387 ); 
   nand2 U1418 ( L2536, L2537, L2538 ); 
   nand2 U1419 ( L3272, L3275, L2539 ); 
   inv U1420 ( L3334, L3338 ); 
   inv U1421 ( L3342, L3346 ); 
   nand2 U1422 ( L3350, L3353, L2556 ); 
   nand2 U1423 ( L2579, L2580, L2581 ); 
   nand2 U1424 ( L3398, L3401, L2601 ); 
   nand2 U1425 ( L2615, L2616, L2617 ); 
   nand2 U1426 ( L2621, L2622, L2623 ); 
   buffer U1427 ( L2635, L2638 ); 
   inv U1428 ( L3454, L3458 ); 
   or3 U1429 ( L2805, L2808, L2811, L2814 ); 
   nor3 U1430 ( L2805, L2808, L2811, L2816 ); 
   nand2 U1431 ( L3264, L3267, L3111 ); 
   nand2 U1432 ( L2539, L2540, L2541 ); 
   nand2 U1433 ( L2556, L2557, L2558 ); 
   inv U1434 ( L3355, L3361 ); 
   nand2 U1435 ( L3355, L3362, L2571 ); 
   inv U1436 ( L3363, L3369 ); 
   nand2 U1437 ( L3363, L3370, L2577 ); 
   inv U1438 ( L3379, L3385 ); 
   nand2 U1439 ( L3379, L3386, L2593 ); 
   inv U1440 ( L3387, L3393 ); 
   nand2 U1441 ( L3387, L3394, L2598 ); 
   nand2 U1442 ( L2601, L2602, L2603 ); 
   nand2 U1443 ( L3111, L3112, L3113 ); 
   and2 U1444 ( L330, L2538, L3116 ); 
   inv U1445 ( L2623, L3451 ); 
   inv U1446 ( L2816, L395 ); 
   nand2 U1447 ( L3358, L3361, L2570 ); 
   nand2 U1448 ( L3366, L3369, L2576 ); 
   nand2 U1449 ( L3382, L3385, L2592 ); 
   nand2 U1450 ( L3390, L3393, L2597 ); 
   and2 U1451 ( L2581, L2733, L2736 ); 
   and2 U1452 ( L2581, L2734, L2739 ); 
   and2 U1453 ( L2617, L2785, L2788 ); 
   buffer U1454 ( L2638, L3438 ); 
   and2 U1455 ( L2617, L2647, L3446 ); 
   buffer U1456 ( L2814, L3459 ); 
   and2 U1457 ( L2814, L395, L396 ); 
   inv U1458 ( L3113, L3119 ); 
   inv U1459 ( L3116, L3120 ); 
   nand2 U1460 ( L2570, L2571, L2572 ); 
   nand2 U1461 ( L2576, L2577, L2578 ); 
   nand2 U1462 ( L2592, L2593, L2594 ); 
   nand2 U1463 ( L2597, L2598, L2599 ); 
   nand2 U1464 ( L3451, L3458, L2677 ); 
   inv U1465 ( L3451, L3457 ); 
   and2 U1466 ( L2558, L2697, L2700 ); 
   and2 U1467 ( L2603, L2768, L2771 ); 
   buffer U1468 ( L2541, L3331 ); 
   buffer U1469 ( L2541, L3339 ); 
   buffer U1470 ( L2558, L3427 ); 
   buffer U1471 ( L2603, L3443 ); 
   nand2 U1472 ( L3116, L3119, L954 ); 
   nand2 U1473 ( L3113, L3120, L955 ); 
   inv U1474 ( L2599, L2600 ); 
   inv U1475 ( L3438, L3442 ); 
   inv U1476 ( L3446, L3450 ); 
   nand2 U1477 ( L3454, L3457, L2676 ); 
   or3 U1478 ( L2736, L2739, L2742, L2745 ); 
   nor3 U1479 ( L2736, L2739, L2742, L2748 ); 
   inv U1480 ( L3459, L3465 ); 
   inv U1481 ( L2578, L3435 ); 
   nand2 U1482 ( L954, L955, L950 ); 
   inv U1483 ( L3331, L3337 ); 
   nand2 U1484 ( L3331, L3338, L2548 ); 
   inv U1485 ( L3339, L3345 ); 
   nand2 U1486 ( L3339, L3346, L2553 ); 
   nor2 U1487 ( L2600, L2650, L2661 ); 
   and4 U1488 ( L2617, L2603, L2594, L2650, L2662 ); 
   inv U1489 ( L3427, L3433 ); 
   inv U1490 ( L3443, L3449 ); 
   nand2 U1491 ( L3443, L3450, L2672 ); 
   nand2 U1492 ( L2676, L2677, L2674 ); 
   and2 U1493 ( L2572, L2716, L2719 ); 
   and2 U1494 ( L2594, L2751, L2754 ); 
   and2 U1495 ( L2572, L2635, L3430 ); 
   inv U1496 ( L2748, L383 ); 
   and2 U1497 ( L950, L943, L951 ); 
   nand2 U1498 ( L3334, L3337, L2547 ); 
   nand2 U1499 ( L3342, L3345, L2552 ); 
   or2 U1500 ( L2661, L2662, L2663 ); 
   nand2 U1501 ( L3435, L3442, L2670 ); 
   inv U1502 ( L3435, L3441 ); 
   nand2 U1503 ( L3446, L3449, L2671 ); 
   inv U1504 ( L2674, L2675 ); 
   buffer U1505 ( L2745, L3491 ); 
   buffer U1506 ( L2745, L3499 ); 
   and2 U1507 ( L2745, L383, L384 ); 
   nand2 U1508 ( L2547, L2548, L2549 ); 
   nand2 U1509 ( L2552, L2553, L2554 ); 
   nand2 U1510 ( L3430, L3433, L2664 ); 
   inv U1511 ( L3430, L3434 ); 
   nand2 U1512 ( L3438, L3441, L2669 ); 
   nand2 U1513 ( L2671, L2672, L2673 ); 
   and2 U1514 ( L2663, L2752, L2757 ); 
   and2 U1515 ( L2675, L2786, L2791 ); 
   or3 U1516 ( L944, L947, L951, L365 ); 
   nor3 U1517 ( L944, L947, L951, L1031 ); 
   inv U1518 ( L2554, L2555 ); 
   nand2 U1519 ( L3427, L3434, L2665 ); 
   nand2 U1520 ( L2669, L2670, L2667 ); 
   and2 U1521 ( L2673, L2769, L2774 ); 
   inv U1522 ( L3491, L3497 ); 
   inv U1523 ( L3499, L3505 ); 
   inv U1524 ( L1031, L366 ); 
   nor2 U1525 ( L2555, L2638, L2658 ); 
   and4 U1526 ( L2572, L2558, L2549, L2638, L2659 ); 
   nand2 U1527 ( L2664, L2665, L2666 ); 
   inv U1528 ( L2667, L2668 ); 
   and2 U1529 ( L2549, L2678, L2681 ); 
   or3 U1530 ( L2754, L2757, L2760, L2763 ); 
   nor3 U1531 ( L2754, L2757, L2760, L2765 ); 
   or3 U1532 ( L2788, L2791, L2794, L2797 ); 
   nor3 U1533 ( L2788, L2791, L2794, L2799 ); 
   and2 U1534 ( L365, L366, L367 ); 
   or2 U1535 ( L2658, L2659, L2660 ); 
   and2 U1536 ( L2666, L2698, L2703 ); 
   and2 U1537 ( L2668, L2717, L2722 ); 
   or3 U1538 ( L2771, L2774, L2777, L2780 ); 
   nor3 U1539 ( L2771, L2774, L2777, L2782 ); 
   inv U1540 ( L2765, L386 ); 
   inv U1541 ( L2799, L392 ); 
   and2 U1542 ( L2660, L2679, L2684 ); 
   buffer U1543 ( L2797, L3462 ); 
   buffer U1544 ( L2763, L3470 ); 
   and2 U1545 ( L2763, L386, L387 ); 
   inv U1546 ( L2782, L389 ); 
   and2 U1547 ( L2797, L392, L393 ); 
   or3 U1548 ( L2700, L2703, L2706, L2709 ); 
   nor3 U1549 ( L2700, L2703, L2706, L2713 ); 
   or3 U1550 ( L2719, L2722, L2725, L2728 ); 
   nor3 U1551 ( L2719, L2722, L2725, L2730 ); 
   and4 U1552 ( L2816, L2799, L2782, L2765, L2922 ); 
   buffer U1553 ( L2780, L3467 ); 
   and2 U1554 ( L2780, L389, L390 ); 
   or3 U1555 ( L2681, L2684, L2687, L2690 ); 
   nor3 U1556 ( L2681, L2684, L2687, L2694 ); 
   nand2 U1557 ( L3462, L3465, L2821 ); 
   inv U1558 ( L3462, L3466 ); 
   inv U1559 ( L3470, L3474 ); 
   buffer U1560 ( L2709, L378 ); 
   inv U1561 ( L2730, L380 ); 
   nand2 U1562 ( L3459, L3466, L2822 ); 
   inv U1563 ( L3467, L3473 ); 
   nand2 U1564 ( L3467, L3474, L2827 ); 
   buffer U1565 ( L2728, L2839 ); 
   and2 U1566 ( L2709, L2871, L2883 ); 
   buffer U1567 ( L2709, L3507 ); 
   buffer U1568 ( L2690, L375 ); 
   and2 U1569 ( L2728, L380, L381 ); 
   nand2 U1570 ( L2821, L2822, L2823 ); 
   nand2 U1571 ( L3470, L3473, L2826 ); 
   and2 U1572 ( L2871, L2690, L2880 ); 
   and4 U1573 ( L2748, L2730, L2713, L2694, L2925 ); 
   and3 U1574 ( L2713, L2694, L2874, L2928 ); 
   buffer U1575 ( L2690, L3510 ); 
   nand2 U1576 ( L2826, L2827, L2828 ); 
   buffer U1577 ( L2839, L3494 ); 
   buffer U1578 ( L2839, L3502 ); 
   inv U1579 ( L3507, L3513 ); 
   buffer U1580 ( L2883, L3544 ); 
   buffer U1581 ( L2883, L3552 ); 
   and2 U1582 ( L2922, L2925, L406 ); 
   and2 U1583 ( L2922, L2925, L2929 ); 
   buffer U1584 ( L2823, L3475 ); 
   buffer U1585 ( L2823, L3483 ); 
   inv U1586 ( L3510, L3514 ); 
   nand2 U1587 ( L3510, L3513, L3515 ); 
   buffer U1588 ( L2880, L3541 ); 
   buffer U1589 ( L2880, L3549 ); 
   inv U1590 ( L406, L407 ); 
   nor2 U1591 ( L2928, L2929, L2930 ); 
   nand2 U1592 ( L3494, L3497, L2842 ); 
   inv U1593 ( L3494, L3498 ); 
   nand2 U1594 ( L3502, L3505, L2852 ); 
   inv U1595 ( L3502, L3506 ); 
   inv U1596 ( L3544, L3548 ); 
   inv U1597 ( L3552, L3556 ); 
   buffer U1598 ( L2828, L3478 ); 
   buffer U1599 ( L2828, L3486 ); 
   nand2 U1600 ( L3507, L3514, L3516 ); 
   and2 U1601 ( L213, L2930, L408 ); 
   inv U1602 ( L3475, L3481 ); 
   inv U1603 ( L3483, L3489 ); 
   nand2 U1604 ( L3491, L3498, L2843 ); 
   nand2 U1605 ( L3499, L3506, L2853 ); 
   inv U1606 ( L3541, L3547 ); 
   nand2 U1607 ( L3541, L3548, L2887 ); 
   nand2 U1608 ( L3549, L3556, L2896 ); 
   inv U1609 ( L3549, L3555 ); 
   nand2 U1610 ( L3515, L3516, L3520 ); 
   inv U1611 ( L408, L409 ); 
   nand2 U1612 ( L3478, L3481, L2831 ); 
   inv U1613 ( L3478, L3482 ); 
   nand2 U1614 ( L3486, L3489, L2836 ); 
   inv U1615 ( L3486, L3490 ); 
   nand2 U1616 ( L2842, L2843, L2844 ); 
   nand2 U1617 ( L2852, L2853, L2848 ); 
   nand2 U1618 ( L3544, L3547, L2886 ); 
   nand2 U1619 ( L3552, L3555, L2895 ); 
   nand2 U1620 ( L3475, L3482, L2832 ); 
   nand2 U1621 ( L3483, L3490, L2837 ); 
   inv U1622 ( L2848, L2849 ); 
   inv U1623 ( L3520, L3524 ); 
   nand2 U1624 ( L2886, L2887, L2888 ); 
   nand2 U1625 ( L2895, L2896, L2891 ); 
   nand2 U1626 ( L2831, L2832, L2833 ); 
   nand2 U1627 ( L2836, L2837, L2838 ); 
   inv U1628 ( L2891, L2892 ); 
   buffer U1629 ( L2844, L3517 ); 
   and3 U1630 ( L2844, L2888, L2900, L2906 ); 
   and3 U1631 ( L2849, L2888, L2903, L2908 ); 
   inv U1632 ( L2838, L2913 ); 
   inv U1633 ( L3517, L3523 ); 
   nand2 U1634 ( L3517, L3524, L2855 ); 
   and3 U1635 ( L2844, L2892, L2903, L2907 ); 
   and3 U1636 ( L2849, L2892, L2900, L2909 ); 
   buffer U1637 ( L2833, L3525 ); 
   buffer U1638 ( L2833, L3533 ); 
   nand2 U1639 ( L3520, L3523, L2854 ); 
   or4 U1640 ( L2906, L2907, L2908, L2909, L2910 ); 
   buffer U1641 ( L2913, L3560 ); 
   buffer U1642 ( L2913, L3568 ); 
   nand2 U1643 ( L2854, L2855, L2856 ); 
   inv U1644 ( L3533, L3539 ); 
   inv U1645 ( L3525, L3531 ); 
   inv U1646 ( L3568, L3572 ); 
   inv U1647 ( L3560, L3564 ); 
   buffer U1648 ( L2910, L3557 ); 
   buffer U1649 ( L2910, L3565 ); 
   buffer U1650 ( L2856, L3528 ); 
   buffer U1651 ( L2856, L3536 ); 
   nand2 U1652 ( L3557, L3564, L2921 ); 
   nand2 U1653 ( L3565, L3572, L2917 ); 
   inv U1654 ( L3565, L3571 ); 
   inv U1655 ( L3557, L3563 ); 
   nand2 U1656 ( L3528, L3531, L2863 ); 
   nand2 U1657 ( L3536, L3539, L2859 ); 
   nand2 U1658 ( L3560, L3563, L2920 ); 
   nand2 U1659 ( L3568, L3571, L2916 ); 
   inv U1660 ( L3536, L3540 ); 
   inv U1661 ( L3528, L3532 ); 
   nand2 U1662 ( L3525, L3532, L2864 ); 
   nand2 U1663 ( L3533, L3540, L2860 ); 
   nand2 U1664 ( L2920, L2921, L403 ); 
   nand2 U1665 ( L2916, L2917, L404 ); 
   nand2 U1666 ( L2863, L2864, L400 ); 
   nand2 U1667 ( L2859, L2860, L401 ); 
   and2 U1668 ( L403, L404, L405 ); 
   nand2 U1669 ( L400, L401, L402 ); 
endmodule

