// Benchmark "./benchmarks/iscas85/c2670" written by ABC on Sun Apr 28 12:32:38 2024

module c2670  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241,
    G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253,
    G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269,
    G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452, G483,
    G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384,
    G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066,
    G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106,
    G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179,
    G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193,
    G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205,
    G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240,
    G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252,
    G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268,
    G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452,
    G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348,
    G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996,
    G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105,
    G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474,
    G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_G546, new_G560, new_G1385, new_G157, new_G547, new_G258, new_G480,
    new_G486, new_G654, new_G655, new_G658, new_G772, new_G795, new_G865,
    new_G875, new_G882, new_G1251, new_G1254, new_G1261, new_G1284,
    new_G1344, new_G1351, new_G1394, new_G1418, new_G2433, new_G2434,
    new_G2441, new_G2442, new_G2449, new_G2450, new_G2478, new_G1631,
    new_G1655, new_G1710, new_G1721, new_G2682, new_G1955, new_G1959,
    new_G1964, new_G1969, new_G1974, new_G1979, new_G1984, new_G1989,
    new_G1994, new_G1999, new_G2001, new_G2012, new_G2070, new_G2076,
    new_G2082, new_G2088, new_G2094, new_G2099, new_G2103, new_G2457,
    new_G2458, new_G2461, new_G2464, new_G2471, new_G2479, new_G2482,
    new_G2487, new_G2490, new_G2495, new_G2498, new_G2505, new_G2508,
    new_G2675, new_G2683, new_G2686, new_G2691, new_G2694, new_G2699,
    new_G2702, new_G487, new_G1475, new_G1476, new_G1484, new_G1485,
    new_G1493, new_G1494, new_G2459, new_G2460, new_G216, new_G1253,
    new_G1256, new_G558, new_G748, new_G784, new_G807, new_G821, new_G825,
    new_G829, new_G833, new_G837, new_G881, new_G994, new_G1273, new_G1296,
    new_G1310, new_G1314, new_G1318, new_G1322, new_G1326, new_G1406,
    new_G1430, new_G1444, new_G1448, new_G1452, new_G1456, new_G1460,
    new_G1477, new_G1486, new_G1495, new_G2477, new_G1499, new_G2485,
    new_G2486, new_G2493, new_G2494, new_G1643, new_G1667, new_G1681,
    new_G1685, new_G1689, new_G1693, new_G1697, new_G1716, new_G1728,
    new_G2681, new_G1776, new_G2689, new_G2690, new_G2697, new_G2698,
    new_G1831, new_G1893, new_G2007, new_G2018, new_G2467, new_G2468,
    new_G2501, new_G2502, new_G2511, new_G2512, new_G2518, new_G2551,
    new_G2559, new_G2567, new_G2575, new_G2583, new_G2591, new_G2599,
    new_G2607, new_G2615, new_G2623, new_G2705, new_G2706, new_G2735,
    new_G2743, new_G2751, new_G2759, new_G2767, new_G2775, new_G550,
    new_G552, new_G894, new_G1498, new_G1507, new_G1508, new_G1516,
    new_G1517, new_G1775, new_G1784, new_G1785, new_G1793, new_G1794,
    new_G2469, new_G2470, new_G2503, new_G2504, new_G2513, new_G2514,
    new_G2707, new_G2708, new_G551, new_G553, new_G818, new_G819, new_G820,
    new_G822, new_G823, new_G824, new_G826, new_G827, new_G828, new_G830,
    new_G831, new_G832, new_G834, new_G835, new_G836, new_G1307, new_G1308,
    new_G1309, new_G1311, new_G1312, new_G1313, new_G1315, new_G1316,
    new_G1317, new_G1319, new_G1320, new_G1321, new_G1323, new_G1324,
    new_G1325, new_G1441, new_G1442, new_G1443, new_G1445, new_G1446,
    new_G1447, new_G1449, new_G1450, new_G1451, new_G1453, new_G1454,
    new_G1455, new_G1457, new_G1458, new_G1459, new_G1481, new_G1490,
    new_G1500, new_G1509, new_G1518, new_G1521, new_G1525, new_G2557,
    new_G2565, new_G2573, new_G2581, new_G2589, new_G2597, new_G2605,
    new_G2613, new_G2621, new_G2629, new_G1678, new_G1679, new_G1680,
    new_G1682, new_G1683, new_G1684, new_G1686, new_G1687, new_G1688,
    new_G1690, new_G1691, new_G1692, new_G1694, new_G1695, new_G1696,
    new_G1734, new_G1736, new_G1738, new_G1740, new_G1742, new_G1744,
    new_G1746, new_G1748, new_G1750, new_G1777, new_G1786, new_G1795,
    new_G2023, new_G2025, new_G2027, new_G2029, new_G2031, new_G2033,
    new_G2035, new_G2037, new_G2741, new_G2749, new_G2757, new_G2765,
    new_G2773, new_G2781, new_G2515, new_G2522, new_G2525, new_G2528,
    new_G2730, new_G554, new_G838, new_G841, new_G846, new_G854, new_G857,
    new_G1327, new_G1329, new_G1331, new_G1333, new_G1335, new_G1461,
    new_G1464, new_G1467, new_G1470, new_G1473, new_G1698, new_G1701,
    new_G1704, new_G1707, new_G2634, new_G1504, new_G1513, new_G1524,
    new_G1528, new_G1529, new_G1533, new_G1538, new_G1541, new_G1781,
    new_G1790, new_G1806, new_G1810, new_G2734, new_G2521, new_G2524,
    new_G2531, new_G2532, new_G144, new_G147, new_G152, new_G175, new_G187,
    new_G516, new_G852, new_G885, new_G887, new_G893, new_G1028, new_G1031,
    new_G1035, new_G1041, new_G1049, new_G1057, new_G1060, new_G1066,
    new_G1072, new_G1078, new_G1213, new_G1218, new_G1250, new_G1387,
    new_G1389, new_G1537, new_G1540, new_G1735, new_G1737, new_G1739,
    new_G1741, new_G1743, new_G1745, new_G1747, new_G1749, new_G1751,
    new_G2638, new_G2024, new_G2026, new_G2028, new_G2030, new_G2032,
    new_G2034, new_G2036, new_G2038, new_G2154, new_G2523, new_G2533,
    new_G2534, new_G2631, new_G2639, new_G2642, new_G2647, new_G2650,
    new_G2655, new_G2658, new_G2665, new_G2668, new_G1532, new_G1536,
    new_G1539, new_G1542, new_G1544, new_G1547, new_G2065, new_G1809,
    new_G1813, new_G1821, new_G1824, new_G2538, new_G2546, new_G2554,
    new_G2562, new_G2570, new_G2578, new_G2586, new_G2594, new_G2602,
    new_G2610, new_G2618, new_G2626, new_G2738, new_G2746, new_G2754,
    new_G2762, new_G2770, new_G2778, new_G456, new_G466, new_G562,
    new_G883, new_G889, new_G891, new_G1043, new_G1051, new_G1062,
    new_G1068, new_G1074, new_G1080, new_G1225, new_G1227, new_G1232,
    new_G1234, new_G1543, new_G1546, new_G2637, new_G1753, new_G2645,
    new_G2646, new_G2653, new_G2654, new_G1820, new_G1823, new_G2107,
    new_G2110, new_G2118, new_G2123, new_G2151, new_G2158, new_G2161,
    new_G2164, new_G2172, new_G2235, new_G2262, new_G2350, new_G2535,
    new_G2661, new_G2662, new_G2671, new_G2672, new_G468, new_G897,
    new_G898, new_G1228, new_G1235, new_G1545, new_G1548, new_G2542,
    new_G2550, new_G1561, new_G2558, new_G1565, new_G2566, new_G1569,
    new_G2574, new_G1573, new_G2582, new_G1577, new_G2590, new_G1581,
    new_G2598, new_G1585, new_G2606, new_G1589, new_G2614, new_G1593,
    new_G2622, new_G1597, new_G2630, new_G1752, new_G1761, new_G1762,
    new_G1770, new_G1771, new_G1822, new_G1825, new_G2039, new_G2742,
    new_G2043, new_G2750, new_G2047, new_G2758, new_G2051, new_G2766,
    new_G2055, new_G2774, new_G2059, new_G2782, new_G2663, new_G2664,
    new_G2673, new_G2674, new_G146, new_G462, new_G2113, new_G2114,
    new_G2122, new_G2129, new_G592, new_G2167, new_G2168, new_G2176,
    new_G2241, new_G2266, new_G743, new_G749, new_G886, new_G995,
    new_G1006, new_G1550, new_G2354, new_G2541, new_G1562, new_G1566,
    new_G1570, new_G1574, new_G1578, new_G1582, new_G1586, new_G1590,
    new_G1594, new_G1598, new_G1754, new_G1763, new_G1772, new_G2040,
    new_G2044, new_G2048, new_G2052, new_G2056, new_G2060, new_G2115,
    new_G2126, new_G2131, new_G2134, new_G2141, new_G2144, new_G2157,
    new_G2160, new_G2169, new_G2177, new_G2180, new_G2187, new_G2190,
    new_G2207, new_G2254, new_G2334, new_G2342, new_G2422, new_G2543,
    new_G2709, new_G2712, new_G2727, new_G569, new_G570, new_G599,
    new_G600, new_G896, new_G1549, new_G1243, new_G1245, new_G1257,
    new_G1258, new_G1563, new_G1567, new_G1571, new_G1575, new_G1579,
    new_G1583, new_G1587, new_G1591, new_G1595, new_G1599, new_G2041,
    new_G2045, new_G2049, new_G2053, new_G2057, new_G2061, new_G2159,
    new_G475, new_G490, new_G496, new_G502, new_G508, new_G765, new_G769,
    new_G571, new_G2121, new_G579, new_G587, new_G2130, new_G596, new_G601,
    new_G2175, new_G609, new_G2258, new_G1014, new_G1018, new_G717,
    new_G723, new_G729, new_G735, new_G753, new_G2338, new_G999, new_G1091,
    new_G2346, new_G2426, new_G1337, new_G2549, new_G1552, new_G1600,
    new_G1596, new_G1592, new_G1588, new_G1584, new_G1580, new_G1576,
    new_G1572, new_G1568, new_G1564, new_G2062, new_G2058, new_G2054,
    new_G2050, new_G2046, new_G2042, new_G1758, new_G1767, new_G1798,
    new_G1802, new_G2733, new_G1829, new_G2137, new_G2138, new_G2147,
    new_G2148, new_G2183, new_G2184, new_G2193, new_G2194, new_G2210,
    new_G2213, new_G2715, new_G2716, new_G1094, new_G1096, new_G578,
    new_G588, new_G608, new_G742, new_G1005, new_G1092, new_G1551,
    new_G1554, new_G1555, new_G1557, new_G1558, new_G1828, new_G1845,
    new_G1907, new_G2139, new_G2140, new_G2149, new_G2150, new_G2185,
    new_G2186, new_G2195, new_G2196, new_G2717, new_G2718, new_G154,
    new_G155, new_G763, new_G767, new_G531, new_G537, new_G575, new_G580,
    new_G589, new_G605, new_G610, new_G1012, new_G1016, new_G705, new_G711,
    new_G1093, new_G1355, new_G1553, new_G1556, new_G1559, new_G1601,
    new_G1801, new_G1805, new_G1815, new_G1818, new_G1830, new_G1836,
    new_G1850, new_G1898, new_G1912, new_G2197, new_G2200, new_G2214,
    new_G2215, new_G2217, new_G2220, new_G2722, new_G492, new_G498,
    new_G504, new_G510, new_G519, new_G525, new_G533, new_G539, new_G693,
    new_G699, new_G707, new_G713, new_G719, new_G725, new_G731, new_G737,
    new_G1560, new_G1814, new_G1817, new_G2216, new_G493, new_G499,
    new_G505, new_G511, new_G521, new_G527, new_G534, new_G540, new_G584,
    new_G613, new_G617, new_G621, new_G625, new_G676, new_G695, new_G701,
    new_G708, new_G714, new_G720, new_G726, new_G732, new_G738, new_G1087,
    new_G1108, new_G1361, new_G1369, new_G1373, new_G1377, new_G1607,
    new_G1615, new_G1619, new_G1623, new_G1816, new_G1819, new_G2726,
    new_G1842, new_G1858, new_G1863, new_G1866, new_G1868, new_G1870,
    new_G1872, new_G1874, new_G1876, new_G1904, new_G1920, new_G1925,
    new_G1928, new_G1930, new_G1932, new_G1934, new_G1936, new_G1938,
    new_G2203, new_G2204, new_G2223, new_G2224, new_G2238, new_G522,
    new_G528, new_G696, new_G702, new_G1881, new_G1883, new_G1885,
    new_G1887, new_G1889, new_G1891, new_G1943, new_G1945, new_G1947,
    new_G1949, new_G1951, new_G1953, new_G2205, new_G2206, new_G2225,
    new_G2226, new_G2719, new_G616, new_G620, new_G624, new_G628, new_G630,
    new_G633, new_G636, new_G639, new_G645, new_G2242, new_G675, new_G1107,
    new_G1368, new_G1371, new_G1375, new_G1614, new_G1617, new_G1621,
    new_G1856, new_G1861, new_G1918, new_G1923, new_G2230, new_G2246,
    new_G2270, new_G2278, new_G2286, new_G2294, new_G2302, new_G2310,
    new_G2358, new_G2366, new_G2374, new_G2382, new_G2390, new_G2398,
    new_G629, new_G632, new_G635, new_G638, new_G646, new_G677, new_G1827,
    new_G907, new_G915, new_G922, new_G924, new_G937, new_G946, new_G1109,
    new_G1125, new_G1133, new_G1140, new_G1142, new_G1155, new_G1164,
    new_G1378, new_G1380, new_G1382, new_G1624, new_G1626, new_G1628,
    new_G2725, new_G1859, new_G1864, new_G1921, new_G1926, new_G2267,
    new_G2275, new_G2283, new_G2291, new_G2299, new_G2307, new_G2318,
    new_G2326, new_G2355, new_G2363, new_G2371, new_G2379, new_G2387,
    new_G2395, new_G2406, new_G2414, new_G647, new_G631, new_G634,
    new_G637, new_G640, new_G2234, new_G2250, new_G679, new_G1826,
    new_G2274, new_G2282, new_G2290, new_G2298, new_G2306, new_G2314,
    new_G1110, new_G2362, new_G2370, new_G2378, new_G2386, new_G2394,
    new_G2402, new_G1877, new_G1879, new_G1939, new_G1941, new_G143,
    new_G671, new_G674, new_G686, new_G2273, new_G900, new_G2281, new_G909,
    new_G2289, new_G917, new_G2297, new_G926, new_G2305, new_G929,
    new_G2313, new_G939, new_G2322, new_G2330, new_G967, new_G1104,
    new_G1106, new_G2361, new_G1118, new_G2369, new_G1127, new_G2377,
    new_G1135, new_G2385, new_G1144, new_G2393, new_G1147, new_G2401,
    new_G1157, new_G2410, new_G2418, new_G1184, new_G2227, new_G2243,
    new_G2251, new_G2259, new_G2331, new_G2339, new_G2347, new_G2419,
    new_G687, new_G899, new_G908, new_G916, new_G925, new_G928, new_G938,
    new_G954, new_G961, new_G1117, new_G1126, new_G1134, new_G1143,
    new_G1146, new_G1156, new_G1172, new_G1179, new_G2315, new_G2323,
    new_G2403, new_G2411, new_G2233, new_G642, new_G2249, new_G649,
    new_G2257, new_G665, new_G684, new_G2265, new_G688, new_G901, new_G910,
    new_G918, new_G927, new_G930, new_G940, new_G2337, new_G963, new_G2345,
    new_G1099, new_G1115, new_G2353, new_G1119, new_G1128, new_G1136,
    new_G1145, new_G1148, new_G1158, new_G2425, new_G1181, new_G641,
    new_G648, new_G664, new_G683, new_G2321, new_G948, new_G2329, new_G956,
    new_G962, new_G1098, new_G1114, new_G2409, new_G1166, new_G2417,
    new_G1174, new_G1180, new_G643, new_G650, new_G666, new_G681, new_G690,
    new_G947, new_G955, new_G964, new_G968, new_G970, new_G971, new_G972,
    new_G978, new_G979, new_G1100, new_G1112, new_G1165, new_G1173,
    new_G1182, new_G1185, new_G1187, new_G1188, new_G1189, new_G1195,
    new_G1196, new_G644, new_G884, new_G949, new_G957, new_G969, new_G973,
    new_G1167, new_G1175, new_G1186, new_G1190, new_G680, new_G682,
    new_G895, new_G1025, new_G1111, new_G1113, new_G685, new_G976,
    new_G977, new_G980, new_G981, new_G1116, new_G1193, new_G1194,
    new_G1197, new_G1198, new_G982, new_G983, new_G988, new_G1027,
    new_G1199, new_G1200, new_G1205, new_G984, new_G1085, new_G1201,
    new_G987, new_G990, new_G1204, new_G1207, new_G989, new_G1206,
    new_G991, new_G1208, new_G1221, new_G1238, new_G1239, new_G1240,
    new_G1247, new_G471, new_G473, new_G1088, new_G1089;
  assign G350 = G452;
  assign G335 = G452;
  assign G409 = G452;
  assign new_G546 = G1 & G3;
  assign new_G560 = ~G559;
  assign G369 = G1083;
  assign G367 = G1083;
  assign new_G1385 = ~G1384;
  assign G411 = G2066;
  assign G337 = G2066;
  assign G384 = G2066;
  assign new_G157 = G2072 & G2078 & G2090 & G2084;
  assign new_G547 = ~new_G546;
  assign G218 = ~G44;
  assign G219 = ~G132;
  assign G220 = ~G82;
  assign G221 = ~G96;
  assign G235 = ~G69;
  assign G236 = ~G120;
  assign G237 = ~G57;
  assign G238 = ~G108;
  assign new_G258 = G661 & G2 & G15;
  assign new_G480 = G661;
  assign new_G486 = G37 & G37;
  assign new_G654 = G452;
  assign new_G655 = G8;
  assign new_G658 = G8;
  assign new_G772 = G543;
  assign new_G795 = G651;
  assign new_G865 = ~G860;
  assign new_G875 = ~G868;
  assign new_G882 = G11 & G868;
  assign new_G1251 = G44 & G96 & G132 & G82;
  assign new_G1254 = G69 & G108 & G120 & G57;
  assign new_G1261 = G543;
  assign new_G1284 = G651;
  assign new_G1344 = ~G1341;
  assign new_G1351 = ~G1348;
  assign new_G1394 = G2104;
  assign new_G1418 = G2105;
  assign new_G2433 = ~G2427;
  assign new_G2434 = ~G2430;
  assign new_G2441 = ~G2435;
  assign new_G2442 = ~G2438;
  assign new_G2449 = ~G2443;
  assign new_G2450 = ~G2446;
  assign new_G2478 = ~G2474;
  assign new_G1631 = G2104;
  assign new_G1655 = G2105;
  assign new_G1710 = G16;
  assign new_G1721 = G16;
  assign new_G2682 = ~G2678;
  assign new_G1955 = G7 & G661;
  assign new_G1959 = ~G1956;
  assign new_G1964 = ~G1961;
  assign new_G1969 = ~G1966;
  assign new_G1974 = ~G1971;
  assign new_G1979 = ~G1976;
  assign new_G1984 = ~G1981;
  assign new_G1989 = ~G1986;
  assign new_G1994 = ~G1991;
  assign new_G1999 = ~G1996;
  assign new_G2001 = G29;
  assign new_G2012 = G29;
  assign new_G2070 = ~G2067;
  assign new_G2076 = ~G2072;
  assign new_G2082 = ~G2078;
  assign new_G2088 = ~G2084;
  assign new_G2094 = ~G2090;
  assign new_G2099 = ~G2096;
  assign new_G2103 = ~G2100;
  assign new_G2457 = ~G2451;
  assign new_G2458 = ~G2454;
  assign new_G2461 = G1348;
  assign new_G2464 = G1341;
  assign new_G2471 = G1956;
  assign new_G2479 = G1966;
  assign new_G2482 = G1961;
  assign new_G2487 = G1976;
  assign new_G2490 = G1971;
  assign new_G2495 = G1986;
  assign new_G2498 = G1981;
  assign new_G2505 = G1996;
  assign new_G2508 = G1991;
  assign new_G2675 = G2067;
  assign new_G2683 = G2078;
  assign new_G2686 = G2072;
  assign new_G2691 = G2090;
  assign new_G2694 = G2084;
  assign new_G2699 = G2100;
  assign new_G2702 = G2096;
  assign G158 = ~new_G157;
  assign G259 = ~new_G258;
  assign new_G487 = ~new_G486;
  assign G391 = new_G654;
  assign new_G1475 = ~G2430 | ~new_G2433;
  assign new_G1476 = ~G2427 | ~new_G2434;
  assign new_G1484 = ~G2438 | ~new_G2441;
  assign new_G1485 = ~G2435 | ~new_G2442;
  assign new_G1493 = ~G2446 | ~new_G2449;
  assign new_G1494 = ~G2443 | ~new_G2450;
  assign new_G2459 = ~G2454 | ~new_G2457;
  assign new_G2460 = ~G2451 | ~new_G2458;
  assign G173 = G94 & new_G654;
  assign new_G216 = G2106 & new_G1955;
  assign G223 = ~new_G1955;
  assign G234 = ~G567 | ~new_G1955;
  assign new_G1253 = ~new_G1251;
  assign new_G1256 = ~new_G1254;
  assign new_G558 = new_G1254 & new_G1251;
  assign new_G748 = new_G655;
  assign new_G784 = ~new_G772;
  assign new_G807 = ~new_G795;
  assign new_G821 = new_G795 & G80 & new_G772;
  assign new_G825 = new_G795 & G68 & new_G772;
  assign new_G829 = new_G795 & G79 & new_G772;
  assign new_G833 = new_G795 & G78 & new_G772;
  assign new_G837 = new_G795 & G77 & new_G772;
  assign new_G881 = G11 & new_G875;
  assign new_G994 = new_G655;
  assign new_G1273 = ~new_G1261;
  assign new_G1296 = ~new_G1284;
  assign new_G1310 = new_G1284 & G76 & new_G1261;
  assign new_G1314 = new_G1284 & G75 & new_G1261;
  assign new_G1318 = new_G1284 & G74 & new_G1261;
  assign new_G1322 = new_G1284 & G73 & new_G1261;
  assign new_G1326 = new_G1284 & G72 & new_G1261;
  assign new_G1406 = ~new_G1394;
  assign new_G1430 = ~new_G1418;
  assign new_G1444 = new_G1418 & G114 & new_G1394;
  assign new_G1448 = new_G1418 & G113 & new_G1394;
  assign new_G1452 = new_G1418 & G112 & new_G1394;
  assign new_G1456 = new_G1418 & G111 & new_G1394;
  assign new_G1460 = new_G1394 & new_G1418;
  assign new_G1477 = ~new_G1475 | ~new_G1476;
  assign new_G1486 = ~new_G1484 | ~new_G1485;
  assign new_G1495 = ~new_G1493 | ~new_G1494;
  assign new_G2477 = ~new_G2471;
  assign new_G1499 = ~new_G2471 | ~new_G2478;
  assign new_G2485 = ~new_G2479;
  assign new_G2486 = ~new_G2482;
  assign new_G2493 = ~new_G2487;
  assign new_G2494 = ~new_G2490;
  assign new_G1643 = ~new_G1631;
  assign new_G1667 = ~new_G1655;
  assign new_G1681 = new_G1655 & G118 & new_G1631;
  assign new_G1685 = new_G1655 & G107 & new_G1631;
  assign new_G1689 = new_G1655 & G117 & new_G1631;
  assign new_G1693 = new_G1655 & G116 & new_G1631;
  assign new_G1697 = new_G1655 & G115 & new_G1631;
  assign new_G1716 = ~new_G1710;
  assign new_G1728 = ~new_G1721;
  assign new_G2681 = ~new_G2675;
  assign new_G1776 = ~new_G2675 | ~new_G2682;
  assign new_G2689 = ~new_G2683;
  assign new_G2690 = ~new_G2686;
  assign new_G2697 = ~new_G2691;
  assign new_G2698 = ~new_G2694;
  assign new_G1831 = new_G658;
  assign new_G1893 = new_G658;
  assign new_G2007 = ~new_G2001;
  assign new_G2018 = ~new_G2012;
  assign new_G2467 = ~new_G2461;
  assign new_G2468 = ~new_G2464;
  assign new_G2501 = ~new_G2495;
  assign new_G2502 = ~new_G2498;
  assign new_G2511 = ~new_G2505;
  assign new_G2512 = ~new_G2508;
  assign new_G2518 = ~new_G2459 | ~new_G2460;
  assign new_G2551 = new_G1344;
  assign new_G2559 = new_G1351;
  assign new_G2567 = new_G1959;
  assign new_G2575 = new_G1964;
  assign new_G2583 = new_G1969;
  assign new_G2591 = new_G1974;
  assign new_G2599 = new_G1979;
  assign new_G2607 = new_G1984;
  assign new_G2615 = new_G1989;
  assign new_G2623 = new_G1994;
  assign new_G2705 = ~new_G2699;
  assign new_G2706 = ~new_G2702;
  assign new_G2735 = new_G1999;
  assign new_G2743 = new_G2070;
  assign new_G2751 = new_G2076;
  assign new_G2759 = new_G2082;
  assign new_G2767 = new_G2088;
  assign new_G2775 = new_G2094;
  assign G217 = ~new_G216;
  assign new_G550 = G2106 & new_G1253;
  assign new_G552 = G567 & new_G1256;
  assign G325 = new_G558;
  assign new_G894 = new_G881 | new_G882;
  assign new_G1498 = ~G2474 | ~new_G2477;
  assign new_G1507 = ~new_G2482 | ~new_G2485;
  assign new_G1508 = ~new_G2479 | ~new_G2486;
  assign new_G1516 = ~new_G2490 | ~new_G2493;
  assign new_G1517 = ~new_G2487 | ~new_G2494;
  assign new_G1775 = ~G2678 | ~new_G2681;
  assign new_G1784 = ~new_G2686 | ~new_G2689;
  assign new_G1785 = ~new_G2683 | ~new_G2690;
  assign new_G1793 = ~new_G2694 | ~new_G2697;
  assign new_G1794 = ~new_G2691 | ~new_G2698;
  assign new_G2469 = ~new_G2464 | ~new_G2467;
  assign new_G2470 = ~new_G2461 | ~new_G2468;
  assign new_G2503 = ~new_G2498 | ~new_G2501;
  assign new_G2504 = ~new_G2495 | ~new_G2502;
  assign new_G2513 = ~new_G2508 | ~new_G2511;
  assign new_G2514 = ~new_G2505 | ~new_G2512;
  assign new_G2707 = ~new_G2702 | ~new_G2705;
  assign new_G2708 = ~new_G2699 | ~new_G2706;
  assign G261 = ~new_G558;
  assign new_G551 = ~new_G550;
  assign new_G553 = ~new_G552;
  assign new_G818 = new_G807 & G93 & new_G784;
  assign new_G819 = new_G807 & G55 & new_G772;
  assign new_G820 = new_G795 & G67 & new_G784;
  assign new_G822 = new_G807 & G81 & new_G784;
  assign new_G823 = new_G807 & G43 & new_G772;
  assign new_G824 = new_G795 & G56 & new_G784;
  assign new_G826 = new_G807 & G92 & new_G784;
  assign new_G827 = new_G807 & G54 & new_G772;
  assign new_G828 = new_G795 & G66 & new_G784;
  assign new_G830 = new_G807 & G91 & new_G784;
  assign new_G831 = new_G807 & G53 & new_G772;
  assign new_G832 = new_G795 & G65 & new_G784;
  assign new_G834 = new_G807 & G90 & new_G784;
  assign new_G835 = new_G807 & G52 & new_G772;
  assign new_G836 = new_G795 & G64 & new_G784;
  assign new_G1307 = new_G1296 & G89 & new_G1273;
  assign new_G1308 = new_G1296 & G51 & new_G1261;
  assign new_G1309 = new_G1284 & G63 & new_G1273;
  assign new_G1311 = new_G1296 & G88 & new_G1273;
  assign new_G1312 = new_G1296 & G50 & new_G1261;
  assign new_G1313 = new_G1284 & G62 & new_G1273;
  assign new_G1315 = new_G1296 & G87 & new_G1273;
  assign new_G1316 = new_G1296 & G49 & new_G1261;
  assign new_G1317 = new_G1273 & new_G1284;
  assign new_G1319 = new_G1296 & G86 & new_G1273;
  assign new_G1320 = new_G1296 & G48 & new_G1261;
  assign new_G1321 = new_G1284 & G61 & new_G1273;
  assign new_G1323 = new_G1296 & G85 & new_G1273;
  assign new_G1324 = new_G1296 & G47 & new_G1261;
  assign new_G1325 = new_G1284 & G60 & new_G1273;
  assign new_G1441 = new_G1430 & G138 & new_G1406;
  assign new_G1442 = new_G1430 & G102 & new_G1394;
  assign new_G1443 = new_G1418 & G126 & new_G1406;
  assign new_G1445 = new_G1430 & G137 & new_G1406;
  assign new_G1446 = new_G1430 & G101 & new_G1394;
  assign new_G1447 = new_G1418 & G125 & new_G1406;
  assign new_G1449 = new_G1430 & G136 & new_G1406;
  assign new_G1450 = new_G1430 & G100 & new_G1394;
  assign new_G1451 = new_G1418 & G124 & new_G1406;
  assign new_G1453 = new_G1430 & G135 & new_G1406;
  assign new_G1454 = new_G1430 & G99 & new_G1394;
  assign new_G1455 = new_G1418 & G123 & new_G1406;
  assign new_G1457 = new_G1406 & new_G1430;
  assign new_G1458 = new_G1394 & new_G1430;
  assign new_G1459 = new_G1406 & new_G1418;
  assign new_G1481 = ~new_G1477;
  assign new_G1490 = ~new_G1486;
  assign new_G1500 = ~new_G1498 | ~new_G1499;
  assign new_G1509 = ~new_G1507 | ~new_G1508;
  assign new_G1518 = ~new_G1516 | ~new_G1517;
  assign new_G1521 = new_G1495;
  assign new_G1525 = new_G1495;
  assign new_G2557 = ~new_G2551;
  assign new_G2565 = ~new_G2559;
  assign new_G2573 = ~new_G2567;
  assign new_G2581 = ~new_G2575;
  assign new_G2589 = ~new_G2583;
  assign new_G2597 = ~new_G2591;
  assign new_G2605 = ~new_G2599;
  assign new_G2613 = ~new_G2607;
  assign new_G2621 = ~new_G2615;
  assign new_G2629 = ~new_G2623;
  assign new_G1678 = new_G1667 & G142 & new_G1643;
  assign new_G1679 = new_G1667 & G106 & new_G1631;
  assign new_G1680 = new_G1655 & G130 & new_G1643;
  assign new_G1682 = new_G1667 & G131 & new_G1643;
  assign new_G1683 = new_G1667 & G95 & new_G1631;
  assign new_G1684 = new_G1655 & G119 & new_G1643;
  assign new_G1686 = new_G1667 & G141 & new_G1643;
  assign new_G1687 = new_G1667 & G105 & new_G1631;
  assign new_G1688 = new_G1655 & G129 & new_G1643;
  assign new_G1690 = new_G1667 & G140 & new_G1643;
  assign new_G1691 = new_G1667 & G104 & new_G1631;
  assign new_G1692 = new_G1655 & G128 & new_G1643;
  assign new_G1694 = new_G1667 & G139 & new_G1643;
  assign new_G1695 = new_G1667 & G103 & new_G1631;
  assign new_G1696 = new_G1655 & G127 & new_G1643;
  assign new_G1734 = G19 & new_G1716;
  assign new_G1736 = G4 & new_G1716;
  assign new_G1738 = G20 & new_G1716;
  assign new_G1740 = G5 & new_G1716;
  assign new_G1742 = G21 & new_G1728;
  assign new_G1744 = G22 & new_G1728;
  assign new_G1746 = G23 & new_G1728;
  assign new_G1748 = G6 & new_G1728;
  assign new_G1750 = G24 & new_G1728;
  assign new_G1777 = ~new_G1775 | ~new_G1776;
  assign new_G1786 = ~new_G1784 | ~new_G1785;
  assign new_G1795 = ~new_G1793 | ~new_G1794;
  assign new_G2023 = G25 & new_G2007;
  assign new_G2025 = G32 & new_G2007;
  assign new_G2027 = G26 & new_G2007;
  assign new_G2029 = G33 & new_G2007;
  assign new_G2031 = G27 & new_G2018;
  assign new_G2033 = G34 & new_G2018;
  assign new_G2035 = G35 & new_G2018;
  assign new_G2037 = G28 & new_G2018;
  assign new_G2741 = ~new_G2735;
  assign new_G2749 = ~new_G2743;
  assign new_G2757 = ~new_G2751;
  assign new_G2765 = ~new_G2759;
  assign new_G2773 = ~new_G2767;
  assign new_G2781 = ~new_G2775;
  assign new_G2515 = ~new_G2469 | ~new_G2470;
  assign new_G2522 = ~new_G2518;
  assign new_G2525 = ~new_G2513 | ~new_G2514;
  assign new_G2528 = ~new_G2503 | ~new_G2504;
  assign new_G2730 = ~new_G2707 | ~new_G2708;
  assign new_G554 = new_G551 & new_G553;
  assign new_G838 = new_G821 | new_G820 | new_G818 | new_G819;
  assign new_G841 = new_G825 | new_G824 | new_G822 | new_G823;
  assign new_G846 = new_G829 | new_G828 | new_G826 | new_G827;
  assign new_G854 = new_G833 | new_G832 | new_G830 | new_G831;
  assign new_G857 = new_G837 | new_G836 | new_G834 | new_G835;
  assign new_G1327 = new_G1310 | new_G1309 | new_G1307 | new_G1308;
  assign new_G1329 = new_G1314 | new_G1313 | new_G1311 | new_G1312;
  assign new_G1331 = new_G1318 | new_G1317 | new_G1315 | new_G1316;
  assign new_G1333 = new_G1322 | new_G1321 | new_G1319 | new_G1320;
  assign new_G1335 = new_G1326 | new_G1325 | new_G1323 | new_G1324;
  assign new_G1461 = new_G1444 | new_G1443 | new_G1441 | new_G1442;
  assign new_G1464 = new_G1448 | new_G1447 | new_G1445 | new_G1446;
  assign new_G1467 = new_G1452 | new_G1451 | new_G1449 | new_G1450;
  assign new_G1470 = new_G1456 | new_G1455 | new_G1453 | new_G1454;
  assign new_G1473 = new_G1460 | new_G1459 | new_G1457 | new_G1458;
  assign new_G1698 = new_G1685 | new_G1684 | new_G1682 | new_G1683;
  assign new_G1701 = new_G1689 | new_G1688 | new_G1686 | new_G1687;
  assign new_G1704 = new_G1693 | new_G1692 | new_G1690 | new_G1691;
  assign new_G1707 = new_G1697 | new_G1696 | new_G1694 | new_G1695;
  assign new_G2634 = new_G1681 | new_G1680 | new_G1678 | new_G1679;
  assign G319 = new_G554;
  assign new_G1504 = ~new_G1500;
  assign new_G1513 = ~new_G1509;
  assign new_G1524 = ~new_G1521;
  assign new_G1528 = ~new_G1525;
  assign new_G1529 = new_G1518;
  assign new_G1533 = new_G1518;
  assign new_G1538 = new_G1521 & new_G1486 & new_G1477;
  assign new_G1541 = new_G1525 & new_G1490 & new_G1481;
  assign new_G1781 = ~new_G1777;
  assign new_G1790 = ~new_G1786;
  assign new_G1806 = new_G1795;
  assign new_G1810 = new_G1795;
  assign new_G2734 = ~new_G2730;
  assign new_G2521 = ~new_G2515;
  assign new_G2524 = ~new_G2515 | ~new_G2522;
  assign new_G2531 = ~new_G2525;
  assign new_G2532 = ~new_G2528;
  assign new_G144 = new_G838 & G860;
  assign new_G147 = new_G846 & G860;
  assign new_G152 = new_G841 & G860;
  assign G160 = ~new_G1464;
  assign G162 = ~new_G1467;
  assign G164 = ~new_G1461;
  assign G166 = ~new_G1329;
  assign G168 = ~new_G1327;
  assign G171 = ~new_G857;
  assign new_G175 = new_G554 & G36 & new_G480 & G483;
  assign new_G187 = new_G547 & new_G554 & new_G480 & G483;
  assign new_G516 = new_G838;
  assign new_G852 = ~new_G846;
  assign new_G885 = new_G841 & new_G875;
  assign new_G887 = new_G846 & new_G875;
  assign new_G893 = new_G1327 & G868;
  assign new_G1028 = ~new_G838;
  assign new_G1031 = ~new_G841;
  assign new_G1035 = ~new_G846;
  assign new_G1041 = new_G854;
  assign new_G1049 = new_G857;
  assign new_G1057 = new_G1327;
  assign new_G1060 = new_G1329;
  assign new_G1066 = new_G1331;
  assign new_G1072 = new_G1333;
  assign new_G1078 = new_G1335;
  assign new_G1213 = ~new_G2099 | ~new_G1470;
  assign new_G1218 = ~new_G2103 | ~new_G1473;
  assign new_G1250 = new_G1704;
  assign new_G1387 = new_G1461 & new_G1385;
  assign new_G1389 = ~new_G1464;
  assign new_G1537 = new_G1524 & new_G1481 & new_G1486;
  assign new_G1540 = new_G1528 & new_G1477 & new_G1490;
  assign new_G1735 = new_G841 & new_G1710;
  assign new_G1737 = new_G846 & new_G1710;
  assign new_G1739 = new_G854 & new_G1710;
  assign new_G1741 = new_G857 & new_G1710;
  assign new_G1743 = new_G1327 & new_G1721;
  assign new_G1745 = new_G1329 & new_G1721;
  assign new_G1747 = new_G1331 & new_G1721;
  assign new_G1749 = new_G1333 & new_G1721;
  assign new_G1751 = new_G1335 & new_G1721;
  assign new_G2638 = ~new_G2634;
  assign new_G2024 = new_G1698 & new_G2001;
  assign new_G2026 = new_G1701 & new_G2001;
  assign new_G2028 = new_G1704 & new_G2001;
  assign new_G2030 = new_G1707 & new_G2001;
  assign new_G2032 = new_G1461 & new_G2012;
  assign new_G2034 = new_G1464 & new_G2012;
  assign new_G2036 = new_G1467 & new_G2012;
  assign new_G2038 = new_G1470 & new_G2012;
  assign new_G2154 = new_G841;
  assign new_G2523 = ~new_G2518 | ~new_G2521;
  assign new_G2533 = ~new_G2528 | ~new_G2531;
  assign new_G2534 = ~new_G2525 | ~new_G2532;
  assign new_G2631 = new_G1698;
  assign new_G2639 = new_G1704;
  assign new_G2642 = new_G1701;
  assign new_G2647 = new_G1461;
  assign new_G2650 = new_G1707;
  assign new_G2655 = new_G1467;
  assign new_G2658 = new_G1464;
  assign new_G2665 = new_G1473;
  assign new_G2668 = new_G1470;
  assign G153 = new_G865 | new_G152;
  assign G176 = ~new_G175;
  assign G188 = ~new_G187;
  assign G299 = new_G1041;
  assign G301 = new_G1049;
  assign G286 = new_G1057;
  assign G303 = new_G1060;
  assign G288 = new_G1066;
  assign G305 = new_G1072;
  assign G290 = new_G1078;
  assign new_G1532 = ~new_G1529;
  assign new_G1536 = ~new_G1533;
  assign new_G1539 = ~new_G1537 & ~new_G1538;
  assign new_G1542 = ~new_G1540 & ~new_G1541;
  assign new_G1544 = new_G1529 & new_G1509 & new_G1500;
  assign new_G1547 = new_G1533 & new_G1513 & new_G1504;
  assign new_G2065 = new_G2037 | new_G2038;
  assign new_G1809 = ~new_G1806;
  assign new_G1813 = ~new_G1810;
  assign new_G1821 = new_G1806 & new_G1786 & new_G1777;
  assign new_G1824 = new_G1810 & new_G1790 & new_G1781;
  assign new_G2538 = ~new_G2523 | ~new_G2524;
  assign new_G2546 = ~new_G2533 | ~new_G2534;
  assign new_G2554 = new_G1734 | new_G1735;
  assign new_G2562 = new_G1736 | new_G1737;
  assign new_G2570 = new_G1738 | new_G1739;
  assign new_G2578 = new_G1740 | new_G1741;
  assign new_G2586 = new_G1742 | new_G1743;
  assign new_G2594 = new_G1744 | new_G1745;
  assign new_G2602 = new_G1746 | new_G1747;
  assign new_G2610 = new_G1748 | new_G1749;
  assign new_G2618 = new_G1750 | new_G1751;
  assign new_G2626 = new_G2023 | new_G2024;
  assign new_G2738 = new_G2025 | new_G2026;
  assign new_G2746 = new_G2027 | new_G2028;
  assign new_G2754 = new_G2029 | new_G2030;
  assign new_G2762 = new_G2031 | new_G2032;
  assign new_G2770 = new_G2033 | new_G2034;
  assign new_G2778 = new_G2035 | new_G2036;
  assign new_G456 = G40 & new_G1389 & new_G1387;
  assign new_G466 = ~new_G1387;
  assign new_G562 = ~new_G560 | ~new_G852;
  assign new_G883 = new_G516 & new_G875;
  assign new_G889 = new_G1049 & G868;
  assign new_G891 = new_G1041 & new_G875;
  assign new_G1043 = ~new_G1041;
  assign new_G1051 = ~new_G1049;
  assign new_G1062 = ~new_G1060;
  assign new_G1068 = ~new_G1066;
  assign new_G1074 = ~new_G1072;
  assign new_G1080 = ~new_G1078;
  assign new_G1225 = new_G2099 & new_G1213;
  assign new_G1227 = new_G1213 & new_G1470;
  assign new_G1232 = new_G2103 & new_G1218;
  assign new_G1234 = new_G1218 & new_G1473;
  assign new_G1543 = new_G1532 & new_G1504 & new_G1509;
  assign new_G1546 = new_G1536 & new_G1500 & new_G1513;
  assign new_G2637 = ~new_G2631;
  assign new_G1753 = ~new_G2631 | ~new_G2638;
  assign new_G2645 = ~new_G2639;
  assign new_G2646 = ~new_G2642;
  assign new_G2653 = ~new_G2647;
  assign new_G2654 = ~new_G2650;
  assign new_G1820 = new_G1809 & new_G1781 & new_G1786;
  assign new_G1823 = new_G1813 & new_G1777 & new_G1790;
  assign new_G2107 = new_G1031;
  assign new_G2110 = new_G1028;
  assign new_G2118 = new_G1035;
  assign new_G2123 = ~new_G1057;
  assign new_G2151 = ~new_G852;
  assign new_G2158 = ~new_G2154;
  assign new_G2161 = new_G1031;
  assign new_G2164 = new_G1028;
  assign new_G2172 = new_G1035;
  assign new_G2235 = new_G516;
  assign new_G2262 = new_G1035;
  assign new_G2350 = new_G1035;
  assign new_G2535 = ~new_G1542 | ~new_G1539;
  assign new_G2661 = ~new_G2655;
  assign new_G2662 = ~new_G2658;
  assign new_G2671 = ~new_G2665;
  assign new_G2672 = ~new_G2668;
  assign new_G468 = new_G466 & G40 & new_G1389;
  assign new_G897 = new_G887 | new_G889;
  assign new_G898 = new_G891 | new_G893;
  assign new_G1228 = new_G1225 | new_G1227;
  assign new_G1235 = new_G1232 | new_G1234;
  assign new_G1545 = ~new_G1543 & ~new_G1544;
  assign new_G1548 = ~new_G1546 & ~new_G1547;
  assign new_G2542 = ~new_G2538;
  assign new_G2550 = ~new_G2546;
  assign new_G1561 = ~new_G2554 | ~new_G2557;
  assign new_G2558 = ~new_G2554;
  assign new_G1565 = ~new_G2562 | ~new_G2565;
  assign new_G2566 = ~new_G2562;
  assign new_G1569 = ~new_G2570 | ~new_G2573;
  assign new_G2574 = ~new_G2570;
  assign new_G1573 = ~new_G2578 | ~new_G2581;
  assign new_G2582 = ~new_G2578;
  assign new_G1577 = ~new_G2586 | ~new_G2589;
  assign new_G2590 = ~new_G2586;
  assign new_G1581 = ~new_G2594 | ~new_G2597;
  assign new_G2598 = ~new_G2594;
  assign new_G1585 = ~new_G2602 | ~new_G2605;
  assign new_G2606 = ~new_G2602;
  assign new_G1589 = ~new_G2610 | ~new_G2613;
  assign new_G2614 = ~new_G2610;
  assign new_G1593 = ~new_G2618 | ~new_G2621;
  assign new_G2622 = ~new_G2618;
  assign new_G1597 = ~new_G2626 | ~new_G2629;
  assign new_G2630 = ~new_G2626;
  assign new_G1752 = ~new_G2634 | ~new_G2637;
  assign new_G1761 = ~new_G2642 | ~new_G2645;
  assign new_G1762 = ~new_G2639 | ~new_G2646;
  assign new_G1770 = ~new_G2650 | ~new_G2653;
  assign new_G1771 = ~new_G2647 | ~new_G2654;
  assign new_G1822 = ~new_G1820 & ~new_G1821;
  assign new_G1825 = ~new_G1823 & ~new_G1824;
  assign new_G2039 = ~new_G2738 | ~new_G2741;
  assign new_G2742 = ~new_G2738;
  assign new_G2043 = ~new_G2746 | ~new_G2749;
  assign new_G2750 = ~new_G2746;
  assign new_G2047 = ~new_G2754 | ~new_G2757;
  assign new_G2758 = ~new_G2754;
  assign new_G2051 = ~new_G2762 | ~new_G2765;
  assign new_G2766 = ~new_G2762;
  assign new_G2055 = ~new_G2770 | ~new_G2773;
  assign new_G2774 = ~new_G2770;
  assign new_G2059 = ~new_G2778 | ~new_G2781;
  assign new_G2782 = ~new_G2778;
  assign new_G2663 = ~new_G2658 | ~new_G2661;
  assign new_G2664 = ~new_G2655 | ~new_G2662;
  assign new_G2673 = ~new_G2668 | ~new_G2671;
  assign new_G2674 = ~new_G2665 | ~new_G2672;
  assign new_G146 = new_G562 & new_G865;
  assign new_G462 = ~new_G456;
  assign new_G2113 = ~new_G2107;
  assign new_G2114 = ~new_G2110;
  assign new_G2122 = ~new_G2118;
  assign new_G2129 = ~new_G2123;
  assign new_G592 = new_G562;
  assign new_G2167 = ~new_G2161;
  assign new_G2168 = ~new_G2164;
  assign new_G2176 = ~new_G2172;
  assign new_G2241 = ~new_G2235;
  assign new_G2266 = ~new_G2262;
  assign new_G743 = ~new_G456;
  assign new_G749 = new_G456;
  assign new_G886 = new_G562 & G868;
  assign G284 = new_G897;
  assign G321 = new_G897;
  assign G297 = new_G898;
  assign G280 = new_G898;
  assign new_G995 = new_G456;
  assign new_G1006 = ~new_G456;
  assign new_G1550 = ~new_G2535 | ~new_G2542;
  assign new_G2354 = ~new_G2350;
  assign new_G2541 = ~new_G2535;
  assign new_G1562 = ~new_G2551 | ~new_G2558;
  assign new_G1566 = ~new_G2559 | ~new_G2566;
  assign new_G1570 = ~new_G2567 | ~new_G2574;
  assign new_G1574 = ~new_G2575 | ~new_G2582;
  assign new_G1578 = ~new_G2583 | ~new_G2590;
  assign new_G1582 = ~new_G2591 | ~new_G2598;
  assign new_G1586 = ~new_G2599 | ~new_G2606;
  assign new_G1590 = ~new_G2607 | ~new_G2614;
  assign new_G1594 = ~new_G2615 | ~new_G2622;
  assign new_G1598 = ~new_G2623 | ~new_G2630;
  assign new_G1754 = ~new_G1752 | ~new_G1753;
  assign new_G1763 = ~new_G1761 | ~new_G1762;
  assign new_G1772 = ~new_G1770 | ~new_G1771;
  assign new_G2040 = ~new_G2735 | ~new_G2742;
  assign new_G2044 = ~new_G2743 | ~new_G2750;
  assign new_G2048 = ~new_G2751 | ~new_G2758;
  assign new_G2052 = ~new_G2759 | ~new_G2766;
  assign new_G2056 = ~new_G2767 | ~new_G2774;
  assign new_G2060 = ~new_G2775 | ~new_G2782;
  assign new_G2115 = new_G1043;
  assign new_G2126 = new_G1051;
  assign new_G2131 = new_G1068;
  assign new_G2134 = new_G1062;
  assign new_G2141 = new_G1080;
  assign new_G2144 = new_G1074;
  assign new_G2157 = ~new_G2151;
  assign new_G2160 = ~new_G2151 | ~new_G2158;
  assign new_G2169 = new_G1043;
  assign new_G2177 = new_G1068;
  assign new_G2180 = new_G1062;
  assign new_G2187 = new_G1080;
  assign new_G2190 = new_G1074;
  assign new_G2207 = ~new_G562;
  assign new_G2254 = new_G1043;
  assign new_G2334 = new_G1051;
  assign new_G2342 = new_G1043;
  assign new_G2422 = new_G1051;
  assign new_G2543 = ~new_G1548 | ~new_G1545;
  assign new_G2709 = ~new_G2673 | ~new_G2674;
  assign new_G2712 = ~new_G2663 | ~new_G2664;
  assign new_G2727 = ~new_G1825 | ~new_G1822;
  assign G148 = new_G146 | new_G147;
  assign new_G569 = ~new_G2110 | ~new_G2113;
  assign new_G570 = ~new_G2107 | ~new_G2114;
  assign new_G599 = ~new_G2164 | ~new_G2167;
  assign new_G600 = ~new_G2161 | ~new_G2168;
  assign new_G896 = new_G885 | new_G886;
  assign new_G1549 = ~new_G2538 | ~new_G2541;
  assign new_G1243 = ~new_G1228;
  assign new_G1245 = ~new_G1235;
  assign new_G1257 = new_G468;
  assign new_G1258 = new_G468;
  assign new_G1563 = ~new_G1561 | ~new_G1562;
  assign new_G1567 = ~new_G1565 | ~new_G1566;
  assign new_G1571 = ~new_G1569 | ~new_G1570;
  assign new_G1575 = ~new_G1573 | ~new_G1574;
  assign new_G1579 = ~new_G1577 | ~new_G1578;
  assign new_G1583 = ~new_G1581 | ~new_G1582;
  assign new_G1587 = ~new_G1585 | ~new_G1586;
  assign new_G1591 = ~new_G1589 | ~new_G1590;
  assign new_G1595 = ~new_G1593 | ~new_G1594;
  assign new_G1599 = ~new_G1597 | ~new_G1598;
  assign new_G2041 = ~new_G2039 | ~new_G2040;
  assign new_G2045 = ~new_G2043 | ~new_G2044;
  assign new_G2049 = ~new_G2047 | ~new_G2048;
  assign new_G2053 = ~new_G2051 | ~new_G2052;
  assign new_G2057 = ~new_G2055 | ~new_G2056;
  assign new_G2061 = ~new_G2059 | ~new_G2060;
  assign new_G2159 = ~new_G2154 | ~new_G2157;
  assign new_G475 = new_G462;
  assign new_G490 = new_G1078 & new_G743;
  assign new_G496 = new_G1698 & new_G743;
  assign new_G502 = new_G1701 & new_G743;
  assign new_G508 = new_G1250 & new_G743;
  assign new_G765 = new_G1057 & new_G749;
  assign new_G769 = new_G1060 & new_G749;
  assign new_G571 = ~new_G569 | ~new_G570;
  assign new_G2121 = ~new_G2115;
  assign new_G579 = ~new_G2115 | ~new_G2122;
  assign new_G587 = ~new_G2126 | ~new_G2129;
  assign new_G2130 = ~new_G2126;
  assign new_G596 = ~new_G592;
  assign new_G601 = ~new_G599 | ~new_G600;
  assign new_G2175 = ~new_G2169;
  assign new_G609 = ~new_G2169 | ~new_G2176;
  assign new_G2258 = ~new_G2254;
  assign new_G1014 = new_G1057 & new_G995;
  assign new_G1018 = new_G1060 & new_G995;
  assign new_G717 = new_G1078 & new_G1006;
  assign new_G723 = new_G1698 & new_G1006;
  assign new_G729 = new_G1701 & new_G1006;
  assign new_G735 = new_G1250 & new_G1006;
  assign new_G753 = ~new_G749;
  assign G282 = new_G896;
  assign G323 = new_G896;
  assign new_G2338 = ~new_G2334;
  assign new_G999 = ~new_G995;
  assign new_G1091 = ~new_G1549 | ~new_G1550;
  assign new_G2346 = ~new_G2342;
  assign new_G2426 = ~new_G2422;
  assign new_G1337 = new_G462;
  assign new_G2549 = ~new_G2543;
  assign new_G1552 = ~new_G2543 | ~new_G2550;
  assign new_G1600 = ~new_G1599;
  assign new_G1596 = ~new_G1595;
  assign new_G1592 = ~new_G1591;
  assign new_G1588 = ~new_G1587;
  assign new_G1584 = ~new_G1583;
  assign new_G1580 = ~new_G1579;
  assign new_G1576 = ~new_G1575;
  assign new_G1572 = ~new_G1571;
  assign new_G1568 = ~new_G1567;
  assign new_G1564 = ~new_G1563;
  assign new_G2062 = ~new_G2061;
  assign new_G2058 = ~new_G2057;
  assign new_G2054 = ~new_G2053;
  assign new_G2050 = ~new_G2049;
  assign new_G2046 = ~new_G2045;
  assign new_G2042 = ~new_G2041;
  assign new_G1758 = ~new_G1754;
  assign new_G1767 = ~new_G1763;
  assign new_G1798 = new_G1772;
  assign new_G1802 = new_G1772;
  assign new_G2733 = ~new_G2727;
  assign new_G1829 = ~new_G2727 | ~new_G2734;
  assign new_G2137 = ~new_G2131;
  assign new_G2138 = ~new_G2134;
  assign new_G2147 = ~new_G2141;
  assign new_G2148 = ~new_G2144;
  assign new_G2183 = ~new_G2177;
  assign new_G2184 = ~new_G2180;
  assign new_G2193 = ~new_G2187;
  assign new_G2194 = ~new_G2190;
  assign new_G2210 = ~new_G2159 | ~new_G2160;
  assign new_G2213 = ~new_G2207;
  assign new_G2715 = ~new_G2709;
  assign new_G2716 = ~new_G2712;
  assign new_G1094 = new_G1235 & new_G1245;
  assign new_G1096 = new_G1228 & new_G1243;
  assign new_G578 = ~new_G2118 | ~new_G2121;
  assign new_G588 = ~new_G2123 | ~new_G2130;
  assign new_G608 = ~new_G2172 | ~new_G2175;
  assign new_G742 = new_G1257;
  assign new_G1005 = new_G1257;
  assign new_G1092 = ~new_G1091;
  assign new_G1551 = ~new_G2546 | ~new_G2549;
  assign new_G1554 = new_G1584 & new_G1588 & new_G1592 & new_G1600 & new_G1596;
  assign new_G1555 = new_G1564 & new_G1568 & new_G1572 & new_G1580 & new_G1576;
  assign new_G1557 = new_G2065 & new_G2062;
  assign new_G1558 = new_G2042 & new_G2046 & new_G2050 & new_G2058 & new_G2054;
  assign new_G1828 = ~new_G2730 | ~new_G2733;
  assign new_G1845 = new_G1258;
  assign new_G1907 = new_G1258;
  assign new_G2139 = ~new_G2134 | ~new_G2137;
  assign new_G2140 = ~new_G2131 | ~new_G2138;
  assign new_G2149 = ~new_G2144 | ~new_G2147;
  assign new_G2150 = ~new_G2141 | ~new_G2148;
  assign new_G2185 = ~new_G2180 | ~new_G2183;
  assign new_G2186 = ~new_G2177 | ~new_G2184;
  assign new_G2195 = ~new_G2190 | ~new_G2193;
  assign new_G2196 = ~new_G2187 | ~new_G2194;
  assign new_G2717 = ~new_G2712 | ~new_G2715;
  assign new_G2718 = ~new_G2709 | ~new_G2716;
  assign new_G154 = new_G1094 | new_G1245;
  assign new_G155 = new_G1096 | new_G1243;
  assign new_G763 = new_G1057 & new_G753;
  assign new_G767 = new_G1060 & new_G753;
  assign new_G531 = new_G1066 & new_G753;
  assign new_G537 = new_G1072 & new_G753;
  assign new_G575 = ~new_G571;
  assign new_G580 = ~new_G578 | ~new_G579;
  assign new_G589 = ~new_G587 | ~new_G588;
  assign new_G605 = ~new_G601;
  assign new_G610 = ~new_G608 | ~new_G609;
  assign new_G1012 = new_G1057 & new_G999;
  assign new_G1016 = new_G1060 & new_G999;
  assign new_G705 = new_G1066 & new_G999;
  assign new_G711 = new_G1072 & new_G999;
  assign new_G1093 = new_G1092 & G14;
  assign new_G1355 = new_G475;
  assign new_G1553 = ~new_G1551 | ~new_G1552;
  assign new_G1556 = new_G1554 & new_G1555;
  assign new_G1559 = new_G1557 & new_G1558;
  assign new_G1601 = new_G1337;
  assign new_G1801 = ~new_G1798;
  assign new_G1805 = ~new_G1802;
  assign new_G1815 = new_G1798 & new_G1763 & new_G1754;
  assign new_G1818 = new_G1802 & new_G1767 & new_G1758;
  assign new_G1830 = ~new_G1828 | ~new_G1829;
  assign new_G1836 = new_G475;
  assign new_G1850 = new_G475;
  assign new_G1898 = new_G1337;
  assign new_G1912 = new_G1337;
  assign new_G2197 = ~new_G2149 | ~new_G2150;
  assign new_G2200 = ~new_G2139 | ~new_G2140;
  assign new_G2214 = ~new_G2210;
  assign new_G2215 = ~new_G2210 | ~new_G2213;
  assign new_G2217 = ~new_G2195 | ~new_G2196;
  assign new_G2220 = ~new_G2185 | ~new_G2186;
  assign new_G2722 = ~new_G2717 | ~new_G2718;
  assign G156 = ~new_G154 | ~new_G155;
  assign new_G492 = new_G490 & new_G742;
  assign new_G498 = new_G496 & new_G742;
  assign new_G504 = new_G502 & new_G742;
  assign new_G510 = new_G508 & new_G742;
  assign new_G519 = new_G763 | new_G765;
  assign new_G525 = new_G767 | new_G769;
  assign new_G533 = new_G531 & new_G748;
  assign new_G539 = new_G537 & new_G748;
  assign new_G693 = new_G1012 | new_G1014;
  assign new_G699 = new_G1016 | new_G1018;
  assign new_G707 = new_G705 & new_G994;
  assign new_G713 = new_G711 & new_G994;
  assign new_G719 = new_G717 & new_G1005;
  assign new_G725 = new_G723 & new_G1005;
  assign new_G731 = new_G729 & new_G1005;
  assign new_G737 = new_G735 & new_G1005;
  assign G401 = new_G1093;
  assign new_G1560 = new_G894 & new_G1556 & new_G1559;
  assign new_G1814 = new_G1801 & new_G1758 & new_G1763;
  assign new_G1817 = new_G1805 & new_G1754 & new_G1767;
  assign new_G2216 = ~new_G2207 | ~new_G2214;
  assign G227 = ~new_G1830;
  assign G229 = ~new_G1553;
  assign new_G493 = ~new_G492;
  assign new_G499 = ~new_G498;
  assign new_G505 = ~new_G504;
  assign new_G511 = ~new_G510;
  assign new_G521 = new_G519 & new_G748;
  assign new_G527 = new_G525 & new_G748;
  assign new_G534 = ~new_G533;
  assign new_G540 = ~new_G539;
  assign new_G584 = ~new_G580;
  assign new_G613 = new_G589;
  assign new_G617 = new_G589;
  assign new_G621 = new_G610;
  assign new_G625 = new_G610;
  assign new_G676 = new_G1344 & new_G1355;
  assign new_G695 = new_G693 & new_G994;
  assign new_G701 = new_G699 & new_G994;
  assign new_G708 = ~new_G707;
  assign new_G714 = ~new_G713;
  assign new_G720 = ~new_G719;
  assign new_G726 = ~new_G725;
  assign new_G732 = ~new_G731;
  assign new_G738 = ~new_G737;
  assign new_G1087 = ~new_G1093;
  assign new_G1108 = new_G1344 & new_G1601;
  assign new_G1361 = ~new_G1355;
  assign new_G1369 = new_G1351 & new_G1355;
  assign new_G1373 = new_G1959 & new_G1355;
  assign new_G1377 = new_G1964 & new_G1355;
  assign G311 = new_G1560;
  assign new_G1607 = ~new_G1601;
  assign new_G1615 = new_G1351 & new_G1601;
  assign new_G1619 = new_G1959 & new_G1601;
  assign new_G1623 = new_G1964 & new_G1601;
  assign new_G1816 = ~new_G1814 & ~new_G1815;
  assign new_G1819 = ~new_G1817 & ~new_G1818;
  assign new_G2726 = ~new_G2722;
  assign new_G1842 = ~new_G1836;
  assign new_G1858 = new_G1969 & new_G1836;
  assign new_G1863 = new_G1974 & new_G1836;
  assign new_G1866 = new_G1979 & new_G1836;
  assign new_G1868 = new_G1984 & new_G1836;
  assign new_G1870 = new_G1989 & new_G1850;
  assign new_G1872 = new_G1994 & new_G1850;
  assign new_G1874 = new_G1999 & new_G1850;
  assign new_G1876 = new_G2070 & new_G1850;
  assign new_G1904 = ~new_G1898;
  assign new_G1920 = new_G1969 & new_G1898;
  assign new_G1925 = new_G1974 & new_G1898;
  assign new_G1928 = new_G1979 & new_G1898;
  assign new_G1930 = new_G1984 & new_G1898;
  assign new_G1932 = new_G1989 & new_G1912;
  assign new_G1934 = new_G1994 & new_G1912;
  assign new_G1936 = new_G1999 & new_G1912;
  assign new_G1938 = new_G2070 & new_G1912;
  assign new_G2203 = ~new_G2197;
  assign new_G2204 = ~new_G2200;
  assign new_G2223 = ~new_G2217;
  assign new_G2224 = ~new_G2220;
  assign new_G2238 = ~new_G2215 | ~new_G2216;
  assign G150 = ~new_G1560;
  assign new_G522 = ~new_G521;
  assign new_G528 = ~new_G527;
  assign new_G696 = ~new_G695;
  assign new_G702 = ~new_G701;
  assign new_G1881 = new_G1866 & new_G1831;
  assign new_G1883 = new_G1868 & new_G1831;
  assign new_G1885 = new_G1870 & new_G1845;
  assign new_G1887 = new_G1872 & new_G1845;
  assign new_G1889 = new_G1874 & new_G1845;
  assign new_G1891 = new_G1876 & new_G1845;
  assign new_G1943 = new_G1928 & new_G1893;
  assign new_G1945 = new_G1930 & new_G1893;
  assign new_G1947 = new_G1932 & new_G1907;
  assign new_G1949 = new_G1934 & new_G1907;
  assign new_G1951 = new_G1936 & new_G1907;
  assign new_G1953 = new_G1938 & new_G1907;
  assign new_G2205 = ~new_G2200 | ~new_G2203;
  assign new_G2206 = ~new_G2197 | ~new_G2204;
  assign new_G2225 = ~new_G2220 | ~new_G2223;
  assign new_G2226 = ~new_G2217 | ~new_G2224;
  assign new_G2719 = ~new_G1819 | ~new_G1816;
  assign new_G616 = ~new_G613;
  assign new_G620 = ~new_G617;
  assign new_G624 = ~new_G621;
  assign new_G628 = ~new_G625;
  assign new_G630 = new_G613 & new_G580 & new_G571;
  assign new_G633 = new_G617 & new_G584 & new_G575;
  assign new_G636 = new_G621 & new_G601 & new_G592;
  assign new_G639 = new_G625 & new_G605 & new_G596;
  assign new_G645 = ~new_G2238 | ~new_G2241;
  assign new_G2242 = ~new_G2238;
  assign new_G675 = new_G1999 & new_G1361;
  assign new_G1107 = new_G1999 & new_G1607;
  assign new_G1368 = new_G2070 & new_G1361;
  assign new_G1371 = new_G2076 & new_G1361;
  assign new_G1375 = new_G2082 & new_G1361;
  assign new_G1614 = new_G2070 & new_G1607;
  assign new_G1617 = new_G2076 & new_G1607;
  assign new_G1621 = new_G2082 & new_G1607;
  assign new_G1856 = new_G2088 & new_G1842;
  assign new_G1861 = new_G2094 & new_G1842;
  assign new_G1918 = new_G2088 & new_G1904;
  assign new_G1923 = new_G2094 & new_G1904;
  assign new_G2230 = ~new_G2205 | ~new_G2206;
  assign new_G2246 = ~new_G2225 | ~new_G2226;
  assign new_G2270 = new_G511;
  assign new_G2278 = new_G505;
  assign new_G2286 = new_G499;
  assign new_G2294 = new_G493;
  assign new_G2302 = new_G540;
  assign new_G2310 = new_G534;
  assign new_G2358 = new_G738;
  assign new_G2366 = new_G732;
  assign new_G2374 = new_G726;
  assign new_G2382 = new_G720;
  assign new_G2390 = new_G714;
  assign new_G2398 = new_G708;
  assign new_G629 = new_G616 & new_G575 & new_G580;
  assign new_G632 = new_G620 & new_G571 & new_G584;
  assign new_G635 = new_G624 & new_G596 & new_G601;
  assign new_G638 = new_G628 & new_G592 & new_G605;
  assign new_G646 = ~new_G2235 | ~new_G2242;
  assign new_G677 = new_G675 | new_G676;
  assign new_G1827 = ~new_G2719 | ~new_G2726;
  assign new_G907 = new_G1891 & new_G511;
  assign new_G915 = new_G1889 & new_G505;
  assign new_G922 = new_G1887 & new_G499;
  assign new_G924 = new_G493 & new_G1885;
  assign new_G937 = new_G1883 & new_G540;
  assign new_G946 = new_G1881 & new_G534;
  assign new_G1109 = new_G1107 | new_G1108;
  assign new_G1125 = new_G1953 & new_G738;
  assign new_G1133 = new_G1951 & new_G732;
  assign new_G1140 = new_G1949 & new_G726;
  assign new_G1142 = new_G720 & new_G1947;
  assign new_G1155 = new_G1945 & new_G714;
  assign new_G1164 = new_G1943 & new_G708;
  assign new_G1378 = new_G1368 | new_G1369;
  assign new_G1380 = new_G1371 | new_G1373;
  assign new_G1382 = new_G1375 | new_G1377;
  assign new_G1624 = new_G1614 | new_G1615;
  assign new_G1626 = new_G1617 | new_G1619;
  assign new_G1628 = new_G1621 | new_G1623;
  assign new_G2725 = ~new_G2719;
  assign new_G1859 = new_G1856 | new_G1858;
  assign new_G1864 = new_G1861 | new_G1863;
  assign new_G1921 = new_G1918 | new_G1920;
  assign new_G1926 = new_G1923 | new_G1925;
  assign new_G2267 = new_G1891;
  assign new_G2275 = new_G1889;
  assign new_G2283 = new_G1887;
  assign new_G2291 = new_G1885;
  assign new_G2299 = new_G1883;
  assign new_G2307 = new_G1881;
  assign new_G2318 = new_G528;
  assign new_G2326 = new_G522;
  assign new_G2355 = new_G1953;
  assign new_G2363 = new_G1951;
  assign new_G2371 = new_G1949;
  assign new_G2379 = new_G1947;
  assign new_G2387 = new_G1945;
  assign new_G2395 = new_G1943;
  assign new_G2406 = new_G702;
  assign new_G2414 = new_G696;
  assign new_G647 = ~new_G645 | ~new_G646;
  assign new_G631 = ~new_G629 & ~new_G630;
  assign new_G634 = ~new_G632 & ~new_G633;
  assign new_G637 = ~new_G635 & ~new_G636;
  assign new_G640 = ~new_G638 & ~new_G639;
  assign new_G2234 = ~new_G2230;
  assign new_G2250 = ~new_G2246;
  assign new_G679 = new_G677 & new_G1031;
  assign new_G1826 = ~new_G2722 | ~new_G2725;
  assign new_G2274 = ~new_G2270;
  assign new_G2282 = ~new_G2278;
  assign new_G2290 = ~new_G2286;
  assign new_G2298 = ~new_G2294;
  assign new_G2306 = ~new_G2302;
  assign new_G2314 = ~new_G2310;
  assign new_G1110 = new_G1109 & new_G1031;
  assign new_G2362 = ~new_G2358;
  assign new_G2370 = ~new_G2366;
  assign new_G2378 = ~new_G2374;
  assign new_G2386 = ~new_G2382;
  assign new_G2394 = ~new_G2390;
  assign new_G2402 = ~new_G2398;
  assign new_G1877 = new_G1859 & new_G1831;
  assign new_G1879 = new_G1864 & new_G1831;
  assign new_G1939 = new_G1921 & new_G1893;
  assign new_G1941 = new_G1926 & new_G1893;
  assign new_G143 = new_G647 & new_G865;
  assign new_G671 = new_G1380 & new_G1043;
  assign new_G674 = new_G1378 & new_G1035;
  assign new_G686 = ~new_G1826 | ~new_G1827;
  assign new_G2273 = ~new_G2267;
  assign new_G900 = ~new_G2267 | ~new_G2274;
  assign new_G2281 = ~new_G2275;
  assign new_G909 = ~new_G2275 | ~new_G2282;
  assign new_G2289 = ~new_G2283;
  assign new_G917 = ~new_G2283 | ~new_G2290;
  assign new_G2297 = ~new_G2291;
  assign new_G926 = ~new_G2291 | ~new_G2298;
  assign new_G2305 = ~new_G2299;
  assign new_G929 = ~new_G2299 | ~new_G2306;
  assign new_G2313 = ~new_G2307;
  assign new_G939 = ~new_G2307 | ~new_G2314;
  assign new_G2322 = ~new_G2318;
  assign new_G2330 = ~new_G2326;
  assign new_G967 = new_G1382 & new_G1051;
  assign new_G1104 = new_G1626 & new_G1043;
  assign new_G1106 = new_G1624 & new_G1035;
  assign new_G2361 = ~new_G2355;
  assign new_G1118 = ~new_G2355 | ~new_G2362;
  assign new_G2369 = ~new_G2363;
  assign new_G1127 = ~new_G2363 | ~new_G2370;
  assign new_G2377 = ~new_G2371;
  assign new_G1135 = ~new_G2371 | ~new_G2378;
  assign new_G2385 = ~new_G2379;
  assign new_G1144 = ~new_G2379 | ~new_G2386;
  assign new_G2393 = ~new_G2387;
  assign new_G1147 = ~new_G2387 | ~new_G2394;
  assign new_G2401 = ~new_G2395;
  assign new_G1157 = ~new_G2395 | ~new_G2402;
  assign new_G2410 = ~new_G2406;
  assign new_G2418 = ~new_G2414;
  assign new_G1184 = new_G1628 & new_G1051;
  assign new_G2227 = ~new_G634 | ~new_G631;
  assign new_G2243 = ~new_G640 | ~new_G637;
  assign new_G2251 = new_G1380;
  assign new_G2259 = new_G1378;
  assign new_G2331 = new_G1382;
  assign new_G2339 = new_G1626;
  assign new_G2347 = new_G1624;
  assign new_G2419 = new_G1628;
  assign G145 = new_G143 | new_G144;
  assign new_G687 = ~new_G686;
  assign new_G899 = ~new_G2270 | ~new_G2273;
  assign new_G908 = ~new_G2278 | ~new_G2281;
  assign new_G916 = ~new_G2286 | ~new_G2289;
  assign new_G925 = ~new_G2294 | ~new_G2297;
  assign new_G928 = ~new_G2302 | ~new_G2305;
  assign new_G938 = ~new_G2310 | ~new_G2313;
  assign new_G954 = new_G1879 & new_G528;
  assign new_G961 = new_G1877 & new_G522;
  assign new_G1117 = ~new_G2358 | ~new_G2361;
  assign new_G1126 = ~new_G2366 | ~new_G2369;
  assign new_G1134 = ~new_G2374 | ~new_G2377;
  assign new_G1143 = ~new_G2382 | ~new_G2385;
  assign new_G1146 = ~new_G2390 | ~new_G2393;
  assign new_G1156 = ~new_G2398 | ~new_G2401;
  assign new_G1172 = new_G1941 & new_G702;
  assign new_G1179 = new_G1939 & new_G696;
  assign new_G2315 = new_G1879;
  assign new_G2323 = new_G1877;
  assign new_G2403 = new_G1941;
  assign new_G2411 = new_G1939;
  assign new_G2233 = ~new_G2227;
  assign new_G642 = ~new_G2227 | ~new_G2234;
  assign new_G2249 = ~new_G2243;
  assign new_G649 = ~new_G2243 | ~new_G2250;
  assign new_G2257 = ~new_G2251;
  assign new_G665 = ~new_G2251 | ~new_G2258;
  assign new_G684 = ~new_G2259 | ~new_G2266;
  assign new_G2265 = ~new_G2259;
  assign new_G688 = new_G687 & new_G487;
  assign new_G901 = ~new_G899 | ~new_G900;
  assign new_G910 = ~new_G908 | ~new_G909;
  assign new_G918 = ~new_G916 | ~new_G917;
  assign new_G927 = ~new_G925 | ~new_G926;
  assign new_G930 = ~new_G928 | ~new_G929;
  assign new_G940 = ~new_G938 | ~new_G939;
  assign new_G2337 = ~new_G2331;
  assign new_G963 = ~new_G2331 | ~new_G2338;
  assign new_G2345 = ~new_G2339;
  assign new_G1099 = ~new_G2339 | ~new_G2346;
  assign new_G1115 = ~new_G2347 | ~new_G2354;
  assign new_G2353 = ~new_G2347;
  assign new_G1119 = ~new_G1117 | ~new_G1118;
  assign new_G1128 = ~new_G1126 | ~new_G1127;
  assign new_G1136 = ~new_G1134 | ~new_G1135;
  assign new_G1145 = ~new_G1143 | ~new_G1144;
  assign new_G1148 = ~new_G1146 | ~new_G1147;
  assign new_G1158 = ~new_G1156 | ~new_G1157;
  assign new_G2425 = ~new_G2419;
  assign new_G1181 = ~new_G2419 | ~new_G2426;
  assign new_G641 = ~new_G2230 | ~new_G2233;
  assign new_G648 = ~new_G2246 | ~new_G2249;
  assign new_G664 = ~new_G2254 | ~new_G2257;
  assign new_G683 = ~new_G2262 | ~new_G2265;
  assign G395 = new_G688;
  assign new_G2321 = ~new_G2315;
  assign new_G948 = ~new_G2315 | ~new_G2322;
  assign new_G2329 = ~new_G2323;
  assign new_G956 = ~new_G2323 | ~new_G2330;
  assign new_G962 = ~new_G2334 | ~new_G2337;
  assign new_G1098 = ~new_G2342 | ~new_G2345;
  assign new_G1114 = ~new_G2350 | ~new_G2353;
  assign new_G2409 = ~new_G2403;
  assign new_G1166 = ~new_G2403 | ~new_G2410;
  assign new_G2417 = ~new_G2411;
  assign new_G1174 = ~new_G2411 | ~new_G2418;
  assign new_G1180 = ~new_G2422 | ~new_G2425;
  assign new_G643 = ~new_G641 | ~new_G642;
  assign new_G650 = ~new_G648 | ~new_G649;
  assign new_G666 = ~new_G664 | ~new_G665;
  assign new_G681 = ~new_G683 | ~new_G684;
  assign new_G690 = ~new_G688;
  assign new_G947 = ~new_G2318 | ~new_G2321;
  assign new_G955 = ~new_G2326 | ~new_G2329;
  assign new_G964 = ~new_G962 | ~new_G963;
  assign new_G968 = new_G901 & new_G918 & new_G910 & new_G927;
  assign new_G970 = new_G901 & new_G915;
  assign new_G971 = new_G922 & new_G910 & new_G901;
  assign new_G972 = new_G910 & new_G924 & new_G918 & new_G901;
  assign new_G978 = new_G930 & new_G946;
  assign new_G979 = new_G954 & new_G940 & new_G930;
  assign new_G1100 = ~new_G1098 | ~new_G1099;
  assign new_G1112 = ~new_G1114 | ~new_G1115;
  assign new_G1165 = ~new_G2406 | ~new_G2409;
  assign new_G1173 = ~new_G2414 | ~new_G2417;
  assign new_G1182 = ~new_G1180 | ~new_G1181;
  assign new_G1185 = new_G1119 & new_G1136 & new_G1128 & new_G1145;
  assign new_G1187 = new_G1119 & new_G1133;
  assign new_G1188 = new_G1140 & new_G1128 & new_G1119;
  assign new_G1189 = new_G1128 & new_G1142 & new_G1136 & new_G1119;
  assign new_G1195 = new_G1148 & new_G1164;
  assign new_G1196 = new_G1172 & new_G1158 & new_G1148;
  assign new_G644 = ~new_G643;
  assign new_G884 = new_G650 & G868;
  assign new_G949 = ~new_G947 | ~new_G948;
  assign new_G957 = ~new_G955 | ~new_G956;
  assign new_G969 = ~new_G968;
  assign new_G973 = new_G972 | new_G971 | new_G907 | new_G970;
  assign new_G1167 = ~new_G1165 | ~new_G1166;
  assign new_G1175 = ~new_G1173 | ~new_G1174;
  assign new_G1186 = ~new_G1185;
  assign new_G1190 = new_G1189 | new_G1188 | new_G1125 | new_G1187;
  assign new_G680 = new_G666 & new_G674;
  assign new_G682 = new_G679 & new_G681 & new_G666;
  assign new_G895 = new_G883 | new_G884;
  assign new_G1025 = new_G644 & new_G487;
  assign new_G1111 = new_G1100 & new_G1106;
  assign new_G1113 = new_G1110 & new_G1112 & new_G1100;
  assign new_G685 = new_G682 | new_G671 | new_G680;
  assign G295 = new_G895;
  assign G331 = new_G895;
  assign new_G976 = ~new_G973;
  assign new_G977 = new_G957 & new_G930 & new_G949 & new_G940 & new_G964;
  assign new_G980 = new_G940 & new_G961 & new_G949 & new_G930;
  assign new_G981 = new_G940 & new_G967 & new_G930 & new_G957 & new_G949;
  assign G397 = new_G1025;
  assign new_G1116 = new_G1113 | new_G1104 | new_G1111;
  assign new_G1193 = ~new_G1190;
  assign new_G1194 = new_G1175 & new_G1148 & new_G1167 & new_G1158 & new_G1182;
  assign new_G1197 = new_G1158 & new_G1179 & new_G1167 & new_G1148;
  assign new_G1198 = new_G1158 & new_G1184 & new_G1148 & new_G1175 & new_G1167;
  assign new_G982 = new_G981 | new_G980 | new_G979 | new_G937 | new_G978;
  assign new_G983 = new_G977 & new_G685;
  assign new_G988 = ~new_G976 | ~new_G969;
  assign new_G1027 = ~new_G1025;
  assign new_G1199 = new_G1198 | new_G1197 | new_G1196 | new_G1155 | new_G1195;
  assign new_G1200 = new_G1194 & new_G1116;
  assign new_G1205 = ~new_G1193 | ~new_G1186;
  assign new_G984 = new_G982 | new_G983;
  assign new_G1085 = new_G1830 & new_G690 & new_G1027;
  assign new_G1201 = new_G1199 | new_G1200;
  assign new_G987 = ~new_G984;
  assign new_G990 = new_G988 & new_G984;
  assign new_G1204 = ~new_G1201;
  assign new_G1207 = new_G1205 & new_G1201;
  assign new_G989 = new_G973 & new_G987;
  assign new_G1206 = new_G1190 & new_G1204;
  assign new_G991 = new_G989 | new_G990;
  assign new_G1208 = new_G1206 | new_G1207;
  assign G329 = new_G1208;
  assign new_G1221 = ~new_G1208 | ~new_G991;
  assign new_G1238 = new_G1208 & new_G1221;
  assign new_G1239 = new_G1221 & new_G991;
  assign new_G1240 = new_G1238 | new_G1239;
  assign new_G1247 = ~new_G1240;
  assign new_G471 = new_G1240 & new_G1247;
  assign new_G473 = new_G471 | new_G1247;
  assign G231 = ~new_G473;
  assign new_G1088 = new_G473 & new_G1553 & new_G1087;
  assign new_G1089 = new_G554 & new_G1085 & new_G1088;
  assign G308 = new_G1089;
  assign G225 = ~new_G1089;
endmodule
