// Benchmark "./benchmarks/iscas85/c5315" written by ABC on Sun Apr 28 12:32:39 2024

module c5315  ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_G4114, new_G2825, new_G3547, new_G3549, new_G3551, new_G3553,
    new_G633, new_G814, new_G816, new_G844, new_G846, new_G852, new_G1502,
    new_G1528, new_G1552, new_G1609, new_G1633, new_G1697, new_G1698,
    new_G1701, new_G2179, new_G2203, new_G2226, new_G2281, new_G2304,
    new_G2361, new_G2370, new_G2382, new_G2393, new_G2405, new_G2418,
    new_G2442, new_G2476, new_G2500, new_G2533, new_G2537, new_G2541,
    new_G2545, new_G2549, new_G2553, new_G2557, new_G2561, new_G2627,
    new_G2631, new_G2635, new_G2639, new_G2643, new_G2647, new_G2651,
    new_G2655, new_G2721, new_G2734, new_G2816, new_G2822, new_G2826,
    new_G2828, new_G2882, new_G2886, new_G2890, new_G2894, new_G2898,
    new_G2902, new_G2948, new_G2952, new_G2956, new_G2960, new_G2964,
    new_G2968, new_G3024, new_G3028, new_G3032, new_G3036, new_G3040,
    new_G3044, new_G3048, new_G3052, new_G3092, new_G3105, new_G3175,
    new_G3176, new_G3181, new_G3204, new_G3208, new_G3212, new_G3216,
    new_G3220, new_G3224, new_G3256, new_G3260, new_G3264, new_G3268,
    new_G3272, new_G3276, new_G3302, new_G3314, new_G3354, new_G3358,
    new_G3362, new_G3366, new_G3370, new_G3374, new_G3378, new_G3382,
    new_G3440, new_G3554, new_G3555, new_G3556, new_G3558, new_G3582,
    new_G3616, new_G3628, new_G3660, new_G3684, new_G3721, new_G3728,
    new_G3737, new_G3757, new_G3795, new_G3815, new_G3972, new_G3991,
    new_G4030, new_G4049, new_G4110, new_G4119, new_G4127, new_G4135,
    new_G4143, new_G4151, new_G4159, new_G4167, new_G4175, new_G4183,
    new_G4188, new_G4276, new_G4284, new_G4292, new_G4300, new_G4308,
    new_G4316, new_G4324, new_G4332, new_G4340, new_G4631, new_G4639,
    new_G4647, new_G4655, new_G4663, new_G4671, new_G4676, new_G4764,
    new_G4772, new_G4780, new_G4788, new_G4796, new_G4804, new_G5082,
    new_G5085, new_G5090, new_G5093, new_G5098, new_G5101, new_G5108,
    new_G5111, new_G5332, new_G5335, new_G5340, new_G5343, new_G5348,
    new_G5351, new_G5356, new_G5359, new_G5369, new_G2979, new_G2999,
    new_G1580, new_G1586, new_G1592, new_G1598, new_G1604, new_G1668,
    new_G1674, new_G1680, new_G1686, new_G2254, new_G2260, new_G2266,
    new_G2272, new_G2278, new_G2339, new_G2345, new_G2351, new_G2357,
    new_G711, new_G721, new_G726, new_G731, new_G736, new_G741, new_G746,
    new_G751, new_G756, new_G761, new_G766, new_G771, new_G776, new_G781,
    new_G786, new_G791, new_G796, new_G801, new_G806, new_G3734, new_G842,
    new_G858, new_G881, new_G4123, new_G4131, new_G4139, new_G4147,
    new_G4155, new_G4163, new_G4171, new_G4179, new_G4187, new_G4194,
    new_G4282, new_G4290, new_G4298, new_G4306, new_G4314, new_G4322,
    new_G4330, new_G4338, new_G4346, new_G1526, new_G1540, new_G1564,
    new_G1606, new_G1621, new_G1645, new_G1661, new_G1688, new_G4635,
    new_G4643, new_G4651, new_G4659, new_G4667, new_G4675, new_G4682,
    new_G4770, new_G4778, new_G4786, new_G4794, new_G4802, new_G4810,
    new_G2202, new_G2215, new_G2238, new_G2279, new_G2293, new_G2316,
    new_G2332, new_G2430, new_G2454, new_G2488, new_G2512, new_G2536,
    new_G2540, new_G2544, new_G2548, new_G2552, new_G2556, new_G2560,
    new_G2564, new_G2566, new_G2572, new_G2578, new_G2584, new_G2590,
    new_G2595, new_G2600, new_G2605, new_G2630, new_G2634, new_G2638,
    new_G2642, new_G2646, new_G2650, new_G2654, new_G2658, new_G2660,
    new_G2666, new_G2672, new_G2678, new_G2684, new_G2689, new_G2694,
    new_G2699, new_G2728, new_G2741, new_G2748, new_G2750, new_G2752,
    new_G2754, new_G2756, new_G2758, new_G2760, new_G2762, new_G2764,
    new_G2766, new_G2827, new_G2838, new_G2847, new_G2885, new_G2889,
    new_G2893, new_G2897, new_G2901, new_G2905, new_G2906, new_G2909,
    new_G2913, new_G2918, new_G2922, new_G2927, new_G2951, new_G2955,
    new_G2959, new_G2963, new_G2967, new_G2971, new_G2973, new_G2980,
    new_G2982, new_G2988, new_G2994, new_G3001, new_G3006, new_G3027,
    new_G3031, new_G3035, new_G3039, new_G3043, new_G3047, new_G3051,
    new_G3055, new_G3056, new_G3060, new_G3064, new_G3068, new_G3073,
    new_G3078, new_G3083, new_G3088, new_G3099, new_G3112, new_G3119,
    new_G3121, new_G3123, new_G3125, new_G3126, new_G3128, new_G3130,
    new_G3132, new_G3134, new_G3136, new_G3187, new_G3193, new_G3196,
    new_G3199, new_G3202, new_G3207, new_G3211, new_G3215, new_G3219,
    new_G3223, new_G3227, new_G3228, new_G3232, new_G3234, new_G3238,
    new_G3243, new_G3247, new_G3249, new_G3253, new_G3259, new_G3263,
    new_G3267, new_G3271, new_G3275, new_G3279, new_G3280, new_G3283,
    new_G3287, new_G3292, new_G3295, new_G3299, new_G3305, new_G3306,
    new_G3310, new_G3317, new_G3318, new_G3322, new_G3326, new_G3333,
    new_G3357, new_G3361, new_G3365, new_G3369, new_G3373, new_G3377,
    new_G3381, new_G3385, new_G3386, new_G3390, new_G3394, new_G3398,
    new_G3403, new_G3408, new_G3413, new_G3418, new_G5088, new_G5089,
    new_G5096, new_G5097, new_G3489, new_G3493, new_G3570, new_G3594,
    new_G3622, new_G3632, new_G3637, new_G3640, new_G3643, new_G3646,
    new_G3672, new_G3696, new_G3745, new_G3765, new_G3803, new_G3823,
    new_G5338, new_G5339, new_G5346, new_G5347, new_G5354, new_G5355,
    new_G3979, new_G3998, new_G4037, new_G4056, new_G4094, new_G5104,
    new_G5105, new_G5114, new_G5115, new_G5362, new_G5363, new_G5366,
    new_G5373, new_G2568, new_G2574, new_G2580, new_G2586, new_G2592,
    new_G2597, new_G2602, new_G2607, new_G2662, new_G2668, new_G2674,
    new_G2680, new_G2686, new_G2691, new_G2696, new_G2701, new_G2907,
    new_G2910, new_G2914, new_G2920, new_G2924, new_G2929, new_G2975,
    new_G2984, new_G2990, new_G2996, new_G3003, new_G3008, new_G3015,
    new_G3057, new_G3061, new_G3065, new_G3069, new_G3075, new_G3080,
    new_G3085, new_G3090, new_G3229, new_G3233, new_G3235, new_G3239,
    new_G3244, new_G3250, new_G3254, new_G3281, new_G3284, new_G3288,
    new_G3293, new_G3296, new_G3300, new_G3327, new_G3334, new_G3387,
    new_G3391, new_G3395, new_G3399, new_G3405, new_G3410, new_G3415,
    new_G3420, new_G3422, new_G3423, new_G3431, new_G3432, new_G3895,
    new_G3896, new_G3904, new_G3905, new_G3913, new_G3914, new_G5106,
    new_G5107, new_G5116, new_G5117, new_G5364, new_G5365, new_G2880,
    new_G2881, new_G1579, new_G1585, new_G1591, new_G1597, new_G1603,
    new_G1667, new_G1673, new_G1679, new_G1685, new_G2876, new_G2877,
    new_G2253, new_G2259, new_G2265, new_G2271, new_G2277, new_G2338,
    new_G2344, new_G2350, new_G2356, new_G2868, new_G2869, new_G710,
    new_G2872, new_G2873, new_G720, new_G725, new_G730, new_G735, new_G740,
    new_G745, new_G750, new_G755, new_G760, new_G765, new_G770, new_G775,
    new_G780, new_G785, new_G790, new_G795, new_G800, new_G805, new_G841,
    new_G857, new_G880, new_G1660, new_G2331, new_G2569, new_G2575,
    new_G2581, new_G2587, new_G2593, new_G2598, new_G2603, new_G2608,
    new_G2663, new_G2669, new_G2675, new_G2681, new_G2687, new_G2692,
    new_G2697, new_G2702, new_G2747, new_G2749, new_G2751, new_G2753,
    new_G2755, new_G2757, new_G2759, new_G2761, new_G2763, new_G2765,
    new_G2857, new_G2908, new_G2911, new_G2915, new_G2925, new_G2930,
    new_G2933, new_G2976, new_G2985, new_G2991, new_G2997, new_G3004,
    new_G3009, new_G3058, new_G3062, new_G3066, new_G3070, new_G3076,
    new_G3081, new_G3086, new_G3091, new_G3118, new_G3120, new_G3122,
    new_G3124, new_G3127, new_G3129, new_G3131, new_G3133, new_G3135,
    new_G3147, new_G3192, new_G3195, new_G3198, new_G3201, new_G3230,
    new_G3236, new_G3240, new_G3245, new_G3251, new_G3255, new_G3282,
    new_G3285, new_G3289, new_G3297, new_G3301, new_G3309, new_G3313,
    new_G3321, new_G3325, new_G3328, new_G3329, new_G3335, new_G3336,
    new_G3341, new_G3345, new_G3388, new_G3392, new_G3396, new_G3400,
    new_G3406, new_G3411, new_G3416, new_G3421, new_G3424, new_G3433,
    new_G3492, new_G3496, new_G3780, new_G3783, new_G3786, new_G3789,
    new_G3838, new_G3841, new_G3844, new_G3847, new_G3897, new_G3906,
    new_G3915, new_G4011, new_G4014, new_G4017, new_G4020, new_G4023,
    new_G4069, new_G4072, new_G4075, new_G4078, new_G4081, new_G5206,
    new_G5209, new_G5307, new_G5322, new_G5372, new_G5375, new_G5399,
    new_G2813, new_G3197, new_G3200, new_G3203, new_G3194, new_G2570,
    new_G2576, new_G2582, new_G2588, new_G2664, new_G2670, new_G2676,
    new_G2682, new_G2767, new_G2772, new_G2776, new_G2780, new_G2784,
    new_G2788, new_G2794, new_G2798, new_G2802, new_G2912, new_G2916,
    new_G2936, new_G2977, new_G2986, new_G2992, new_G3059, new_G3063,
    new_G3067, new_G3071, new_G3137, new_G3139, new_G3143, new_G3151,
    new_G3155, new_G3161, new_G3165, new_G3167, new_G3231, new_G3237,
    new_G3241, new_G3286, new_G3290, new_G3330, new_G3337, new_G3342,
    new_G3346, new_G3348, new_G3352, new_G3389, new_G3393, new_G3397,
    new_G3401, new_G3845, new_G5126, new_G5178, new_G5325, new_G5374,
    new_G2810, new_G635, new_G2878, new_G2879, new_G2874, new_G2875,
    new_G703, new_G2866, new_G2867, new_G2870, new_G2871, new_G716,
    new_G819, new_G1789, new_G2036, new_G2611, new_G2615, new_G2619,
    new_G2623, new_G2705, new_G2709, new_G2713, new_G2717, new_G2939,
    new_G2942, new_G2945, new_G3012, new_G3018, new_G3021, new_G3331,
    new_G3338, new_G3343, new_G3347, new_G3428, new_G3437, new_G3514,
    new_G3836, new_G3852, new_G5311, new_G3901, new_G3910, new_G3934,
    new_G3938, new_G4652, new_G4783, new_G5137, new_G5212, new_G5213,
    new_G5260, new_G5263, new_G5268, new_G5271, new_G5276, new_G5279,
    new_G5289, new_G5296, new_G5299, new_G5304, new_G5312, new_G5315,
    new_G5328, new_G5396, new_G5403, new_G1286, new_G2809, new_G597,
    new_G1031, new_G637, new_G671, new_G705, new_G713, new_G1046,
    new_G1064, new_G1071, new_G1097, new_G1111, new_G1128, new_G1145,
    new_G1160, new_G1301, new_G1318, new_G1324, new_G1341, new_G1359,
    new_G1382, new_G1404, new_G1412, new_G1704, new_G1712, new_G1724,
    new_G1742, new_G1749, new_G1775, new_G1806, new_G1823, new_G1829,
    new_G1837, new_G1958, new_G1966, new_G1978, new_G1995, new_G2001,
    new_G2018, new_G2059, new_G2081, new_G2089, new_G2106, new_G3170,
    new_G3332, new_G3339, new_G5132, new_G5184, new_G3853, new_G3874,
    new_G4076, new_G4116, new_G4124, new_G4132, new_G4140, new_G4148,
    new_G4156, new_G4164, new_G4172, new_G4180, new_G4228, new_G4279,
    new_G4287, new_G4295, new_G4303, new_G4311, new_G4319, new_G4327,
    new_G4335, new_G4343, new_G4348, new_G4464, new_G4628, new_G4636,
    new_G4644, new_G4660, new_G4668, new_G4716, new_G4767, new_G4775,
    new_G4791, new_G4799, new_G4807, new_G4812, new_G5118, new_G5121,
    new_G5129, new_G5134, new_G5142, new_G5145, new_G5152, new_G5155,
    new_G5162, new_G5165, new_G5170, new_G5173, new_G5181, new_G5186,
    new_G5189, new_G5196, new_G5199, new_G5214, new_G5215, new_G5329,
    new_G5330, new_G2807, new_G2808, new_G2811, new_G2812, new_G2814,
    new_G2626, new_G2622, new_G2618, new_G2614, new_G2720, new_G2716,
    new_G2712, new_G2708, new_G3731, new_G4658, new_G1777, new_G2019,
    new_G4787, new_G3350, new_G3353, new_G5141, new_G3513, new_G3516,
    new_G3517, new_G3778, new_G3781, new_G3784, new_G3787, new_G3839,
    new_G3842, new_G5266, new_G5267, new_G5274, new_G5275, new_G5302,
    new_G5303, new_G5310, new_G3891, new_G3937, new_G3941, new_G3955,
    new_G3958, new_G4009, new_G4012, new_G4015, new_G4018, new_G4067,
    new_G4070, new_G4073, new_G4079, new_G5239, new_G5282, new_G5283,
    new_G5293, new_G5318, new_G5319, new_G5331, new_G5402, new_G5405,
    new_G595, new_G596, new_G607, new_G608, new_G1845, new_G1846,
    new_G2115, new_G2116, new_G4122, new_G1022, new_G4130, new_G1033,
    new_G4138, new_G1051, new_G4146, new_G1079, new_G4154, new_G1088,
    new_G4162, new_G1099, new_G4170, new_G1115, new_G4178, new_G1133,
    new_G4186, new_G1151, new_G4234, new_G1276, new_G4283, new_G1287,
    new_G4291, new_G1305, new_G4299, new_G1330, new_G4307, new_G1342,
    new_G4315, new_G1363, new_G4323, new_G1388, new_G4331, new_G1420,
    new_G4339, new_G1428, new_G4347, new_G4634, new_G1729, new_G4642,
    new_G1757, new_G4650, new_G1766, new_G1776, new_G4666, new_G1793,
    new_G4674, new_G1811, new_G1849, new_G1852, new_G1875, new_G4722,
    new_G1982, new_G4771, new_G2007, new_G4779, new_G2020, new_G2040,
    new_G4795, new_G2065, new_G4803, new_G2097, new_G4811, new_G2119,
    new_G2122, new_G5124, new_G5125, new_G3452, new_G5133, new_G5140,
    new_G3462, new_G5168, new_G5169, new_G5176, new_G5177, new_G3484,
    new_G5185, new_G3515, new_G3518, new_G3857, new_G3860, new_G3861,
    new_G3869, new_G3870, new_G3878, new_G3881, new_G3882, new_G3890,
    new_G3954, new_G3957, new_G4021, new_G4099, new_G4236, new_G4354,
    new_G4406, new_G4470, new_G4552, new_G4679, new_G4687, new_G4695,
    new_G4703, new_G4711, new_G4724, new_G4818, new_G4855, new_G4865,
    new_G4870, new_G4913, new_G4923, new_G4951, new_G5006, new_G5039,
    new_G5148, new_G5149, new_G5158, new_G5159, new_G5192, new_G5193,
    new_G5202, new_G5203, new_G5284, new_G5285, new_G5320, new_G5321,
    new_G5386, new_G5404, new_G609, new_G1021, new_G1032, new_G1050,
    new_G1078, new_G1087, new_G1098, new_G1114, new_G1132, new_G1150,
    new_G1277, new_G1288, new_G1306, new_G1331, new_G1343, new_G1364,
    new_G1389, new_G1421, new_G1429, new_G1728, new_G1756, new_G1765,
    new_G1778, new_G1792, new_G1810, new_G1983, new_G2008, new_G2021,
    new_G2041, new_G2066, new_G2098, new_G3443, new_G3444, new_G3453,
    new_G3461, new_G3466, new_G3467, new_G3475, new_G3476, new_G3485,
    new_G5243, new_G3862, new_G3871, new_G3883, new_G3892, new_G3956,
    new_G3959, new_G4756, new_G5150, new_G5151, new_G5160, new_G5161,
    new_G5194, new_G5195, new_G5204, new_G5205, new_G5236, new_G5286,
    new_G5379, new_G5389, new_G5425, new_G1023, new_G1034, new_G1052,
    new_G1080, new_G1089, new_G1100, new_G1116, new_G1134, new_G1152,
    new_G4242, new_G1278, new_G1289, new_G1307, new_G1332, new_G1344,
    new_G1365, new_G1390, new_G1422, new_G1430, new_G1730, new_G1758,
    new_G1767, new_G1794, new_G1812, new_G1876, new_G4683, new_G4691,
    new_G4699, new_G4707, new_G4715, new_G4730, new_G1984, new_G2009,
    new_G2042, new_G2067, new_G2099, new_G4869, new_G4927, new_G3445,
    new_G3454, new_G3463, new_G3468, new_G3477, new_G3486, new_G4103,
    new_G4412, new_G4558, new_G4859, new_G4876, new_G4917, new_G4955,
    new_G5012, new_G5043, new_G5216, new_G5219, new_G5226, new_G5229,
    new_G5392, new_G5422, new_G1866, new_G1877, new_G4762, new_G2142,
    new_G2146, new_G5242, new_G3532, new_G3866, new_G3887, new_G3918,
    new_G3922, new_G3926, new_G3930, new_G5429, new_G4104, new_G4743,
    new_G4991, new_G5001, new_G5292, new_G5295, new_G5383, new_G5393,
    new_G5394, new_G1439, new_G1440, new_G1441, new_G1847, new_G1168,
    new_G1169, new_G1170, new_G2117, new_G1086, new_G1166, new_G1171,
    new_G1172, new_G1173, new_G1174, new_G1175, new_G1176, new_G1177,
    new_G1178, new_G1179, new_G1181, new_G1182, new_G1183, new_G1184,
    new_G1188, new_G1189, new_G1190, new_G1191, new_G1192, new_G1193,
    new_G1194, new_G1195, new_G1196, new_G1197, new_G1437, new_G1442,
    new_G1443, new_G1444, new_G1445, new_G1446, new_G1447, new_G1451,
    new_G1454, new_G1455, new_G1456, new_G1457, new_G1465, new_G1466,
    new_G1467, new_G1468, new_G1469, new_G1470, new_G1471, new_G1472,
    new_G1473, new_G1474, new_G1475, new_G1476, new_G1477, new_G1481,
    new_G1482, new_G1764, new_G1843, new_G1850, new_G1851, new_G1853,
    new_G1854, new_G1855, new_G1856, new_G1857, new_G1859, new_G1860,
    new_G1861, new_G1862, new_G1867, new_G1868, new_G1869, new_G1870,
    new_G1871, new_G1872, new_G1873, new_G1874, new_G1878, new_G2113,
    new_G2120, new_G2121, new_G2123, new_G2124, new_G2128, new_G2131,
    new_G2132, new_G2133, new_G2134, new_G2143, new_G2144, new_G2145,
    new_G2147, new_G2148, new_G2149, new_G2150, new_G2151, new_G2152,
    new_G2153, new_G2154, new_G2158, new_G2159, new_G3449, new_G3458,
    new_G3472, new_G3481, new_G3497, new_G3501, new_G3505, new_G3509,
    new_G3531, new_G5428, new_G3967, new_G4191, new_G4199, new_G4207,
    new_G4215, new_G4223, new_G4231, new_G4239, new_G4247, new_G4255,
    new_G4263, new_G4271, new_G4371, new_G4381, new_G4391, new_G4401,
    new_G4429, new_G4439, new_G4449, new_G4459, new_G4497, new_G4507,
    new_G4517, new_G4527, new_G4537, new_G4547, new_G4585, new_G4595,
    new_G4605, new_G4615, new_G4719, new_G4727, new_G4735, new_G4751,
    new_G4759, new_G4835, new_G4845, new_G4893, new_G4903, new_G4961,
    new_G4971, new_G4981, new_G5049, new_G5059, new_G5069, new_G5222,
    new_G5223, new_G5232, new_G5233, new_G5294, new_G5395, new_G589,
    new_G616, new_G619, new_G627, new_G1185, new_G1448, new_G1458,
    new_G1478, new_G1863, new_G4747, new_G2125, new_G2135, new_G2155,
    new_G4995, new_G5005, new_G3533, new_G3921, new_G3925, new_G3929,
    new_G3933, new_G3943, new_G3946, new_G3949, new_G3952, new_G3966,
    new_G4107, new_G4196, new_G4204, new_G4212, new_G4220, new_G4244,
    new_G4252, new_G4260, new_G4268, new_G4361, new_G4419, new_G4467,
    new_G4487, new_G4555, new_G4575, new_G4684, new_G4692, new_G4700,
    new_G4708, new_G4732, new_G4740, new_G4748, new_G4825, new_G4883,
    new_G4928, new_G4941, new_G5009, new_G5029, new_G5224, new_G5225,
    new_G5234, new_G5235, new_G5376, new_G5417, new_G576, new_G1198,
    new_G4195, new_G4203, new_G4211, new_G4219, new_G4227, new_G1217,
    new_G4235, new_G1221, new_G4243, new_G1224, new_G4251, new_G4259,
    new_G4267, new_G4275, new_G1453, new_G4405, new_G4463, new_G4541,
    new_G4551, new_G1895, new_G4723, new_G1899, new_G4731, new_G1902,
    new_G4739, new_G4755, new_G1929, new_G4763, new_G2130, new_G3500,
    new_G3504, new_G3508, new_G3512, new_G3520, new_G3523, new_G3526,
    new_G3529, new_G3837, new_G3942, new_G3945, new_G3948, new_G3951,
    new_G3968, new_G4375, new_G4385, new_G4395, new_G4433, new_G4443,
    new_G4453, new_G4501, new_G4511, new_G4521, new_G4531, new_G4619,
    new_G4589, new_G4599, new_G4609, new_G4839, new_G4849, new_G4897,
    new_G4907, new_G4965, new_G4975, new_G4985, new_G5073, new_G5053,
    new_G5063, new_G5247, new_G5255, new_G590, new_G617, new_G620,
    new_G628, new_G3535, new_G1199, new_G4202, new_G1204, new_G4210,
    new_G1207, new_G4218, new_G1211, new_G4226, new_G1214, new_G1218,
    new_G1222, new_G1225, new_G4250, new_G1237, new_G4258, new_G1242,
    new_G4266, new_G1247, new_G4274, new_G1252, new_G1462, new_G4690,
    new_G1882, new_G4698, new_G1885, new_G4706, new_G1889, new_G4714,
    new_G1892, new_G1896, new_G1900, new_G1903, new_G4738, new_G1915,
    new_G4746, new_G1920, new_G4754, new_G1925, new_G1930, new_G2139,
    new_G3519, new_G3522, new_G3525, new_G3528, new_G3848, new_G3944,
    new_G3947, new_G3950, new_G3953, new_G5421, new_G4111, new_G4112,
    new_G4351, new_G4365, new_G4409, new_G4423, new_G4471, new_G4472,
    new_G4477, new_G4491, new_G4559, new_G4560, new_G4565, new_G4579,
    new_G4815, new_G4829, new_G4873, new_G4887, new_G4931, new_G4934,
    new_G4945, new_G5013, new_G5014, new_G5019, new_G5033, new_G5382,
    new_G5385, new_G3970, new_G1200, new_G1203, new_G1206, new_G1210,
    new_G1213, new_G1219, new_G1223, new_G1236, new_G1241, new_G1246,
    new_G1251, new_G1881, new_G1884, new_G1888, new_G1891, new_G1897,
    new_G1901, new_G1914, new_G1919, new_G1924, new_G1931, new_G3521,
    new_G3524, new_G3527, new_G3530, new_G5251, new_G5259, new_G4113,
    new_G4473, new_G4561, new_G5015, new_G5384, new_G5406, new_G5414,
    new_G1664, new_G2335, new_G718, new_G855, new_G1205, new_G1208,
    new_G1212, new_G1215, new_G1220, new_G1231, new_G1238, new_G1243,
    new_G1248, new_G1253, new_G1272, new_G1483, new_G1883, new_G1886,
    new_G1890, new_G1893, new_G1898, new_G1909, new_G1916, new_G1921,
    new_G1926, new_G1953, new_G2160, new_G4355, new_G4356, new_G4413,
    new_G4414, new_G4474, new_G4481, new_G4562, new_G4569, new_G4819,
    new_G4820, new_G4877, new_G4878, new_G4935, new_G4936, new_G5016,
    new_G5023, new_G5244, new_G5252, new_G5409, new_G566, new_G577,
    new_G3733, new_G1209, new_G1216, new_G1257, new_G1262, new_G1267,
    new_G1887, new_G1894, new_G1935, new_G1943, new_G1948, new_G3779,
    new_G3840, new_G5412, new_G5420, new_G3964, new_G4357, new_G4415,
    new_G4821, new_G4879, new_G4937, new_G567, new_G568, new_G569,
    new_G570, new_G578, new_G579, new_G580, new_G1256, new_G1261,
    new_G1266, new_G1271, new_G1486, new_G1934, new_G1942, new_G1947,
    new_G1952, new_G2163, new_G5250, new_G3537, new_G5258, new_G3542,
    new_G3782, new_G3785, new_G3788, new_G3790, new_G3843, new_G3846,
    new_G3849, new_G3960, new_G5413, new_G3963, new_G4010, new_G4068,
    new_G4358, new_G4416, new_G4480, new_G4483, new_G4568, new_G4571,
    new_G4822, new_G4880, new_G4938, new_G5022, new_G5025, new_G1258,
    new_G1263, new_G1268, new_G1273, new_G1936, new_G1944, new_G1949,
    new_G1954, new_G3536, new_G3541, new_G3791, new_G3792, new_G3793,
    new_G3850, new_G3851, new_G3961, new_G3965, new_G4024, new_G4082,
    new_G4482, new_G4570, new_G5024, new_G1666, new_G1670, new_G2337,
    new_G2341, new_G719, new_G758, new_G798, new_G856, new_G3538,
    new_G3543, new_G3962, new_G4364, new_G4367, new_G4422, new_G4425,
    new_G4484, new_G4572, new_G4828, new_G4831, new_G4886, new_G4889,
    new_G4944, new_G4947, new_G5026, new_G571, new_G572, new_G573,
    new_G574, new_G581, new_G582, new_G583, new_G584, new_G1576, new_G1578,
    new_G659, new_G1672, new_G1676, new_G1678, new_G1682, new_G1684,
    new_G2250, new_G2252, new_G691, new_G2343, new_G2347, new_G2349,
    new_G2353, new_G2355, new_G743, new_G744, new_G748, new_G749, new_G753,
    new_G754, new_G759, new_G783, new_G784, new_G788, new_G789, new_G793,
    new_G794, new_G799, new_G3735, new_G3835, new_G3651, new_G4013,
    new_G4016, new_G4019, new_G4022, new_G4071, new_G4074, new_G4077,
    new_G4080, new_G4096, new_G4366, new_G4424, new_G4830, new_G4888,
    new_G4946, new_G640, new_G662, new_G665, new_G668, new_G674, new_G694,
    new_G697, new_G700, new_G817, new_G839, new_G3540, new_G3545,
    new_G3777, new_G3648, new_G4025, new_G4026, new_G4027, new_G4028,
    new_G4083, new_G4084, new_G4085, new_G4086, new_G4368, new_G4426,
    new_G4490, new_G4493, new_G4578, new_G4581, new_G4832, new_G4890,
    new_G4948, new_G5032, new_G5035, new_G811, new_G812, new_G853,
    new_G878, new_G4492, new_G4580, new_G5034, new_G1582, new_G1584,
    new_G1588, new_G1590, new_G1594, new_G1596, new_G1600, new_G1602,
    new_G2256, new_G2258, new_G2262, new_G2264, new_G2268, new_G2270,
    new_G2274, new_G2276, new_G708, new_G709, new_G723, new_G724, new_G728,
    new_G729, new_G733, new_G734, new_G738, new_G739, new_G768, new_G769,
    new_G773, new_G774, new_G778, new_G779, new_G4374, new_G4377,
    new_G4432, new_G4435, new_G4494, new_G4582, new_G4838, new_G4841,
    new_G4896, new_G4899, new_G4954, new_G4957, new_G5036, new_G643,
    new_G646, new_G649, new_G652, new_G677, new_G680, new_G683, new_G686,
    new_G4376, new_G4434, new_G4840, new_G4898, new_G4956, new_G4378,
    new_G4436, new_G4500, new_G4503, new_G4588, new_G4591, new_G4842,
    new_G4900, new_G4958, new_G5042, new_G5045, new_G4502, new_G4590,
    new_G5044, new_G4384, new_G4387, new_G4442, new_G4445, new_G4504,
    new_G4592, new_G4848, new_G4851, new_G4906, new_G4909, new_G4964,
    new_G4967, new_G5046, new_G4386, new_G4444, new_G4850, new_G4908,
    new_G4966, new_G4388, new_G4446, new_G4510, new_G4513, new_G4598,
    new_G4601, new_G4852, new_G4910, new_G4968, new_G5052, new_G5055,
    new_G4512, new_G4600, new_G5054, new_G4394, new_G4397, new_G4452,
    new_G4455, new_G4514, new_G4602, new_G4858, new_G4861, new_G4916,
    new_G4919, new_G4974, new_G4977, new_G5056, new_G4396, new_G4454,
    new_G4860, new_G4918, new_G4976, new_G4398, new_G4456, new_G4520,
    new_G4523, new_G4608, new_G4611, new_G4862, new_G4920, new_G4978,
    new_G5062, new_G5065, new_G4522, new_G4610, new_G5064, new_G4404,
    new_G1488, new_G4462, new_G1493, new_G4868, new_G2165, new_G4926,
    new_G2170, new_G4524, new_G4612, new_G4984, new_G4987, new_G5066,
    new_G1487, new_G1492, new_G2164, new_G2169, new_G4986, new_G1489,
    new_G1494, new_G2166, new_G2171, new_G4530, new_G4533, new_G4618,
    new_G4543, new_G4988, new_G5072, new_G4997, new_G4532, new_G4542,
    new_G4996, new_G1513, new_G1514, new_G1515, new_G1516, new_G4994,
    new_G2184, new_G2190, new_G2191, new_G2192, new_G2193, new_G4534,
    new_G4544, new_G4998, new_G2183, new_G4620, new_G5074, new_G4540,
    new_G1507, new_G4550, new_G1510, new_G2185, new_G5004, new_G2187,
    new_G1506, new_G1509, new_G4626, new_G2186, new_G2195, new_G5080,
    new_G1508, new_G1511, new_G2188, new_G1512, new_G1518, new_G2189,
    new_G1517, new_G2194, new_G4623, new_G5077, new_G1519, new_G4627,
    new_G2196, new_G5081, new_G1520, new_G2197, new_G1521, new_G2198,
    new_G840, new_G879, new_G1524, new_G2201, new_G3649, new_G3652,
    new_G3657, new_G3658, new_G3636, new_G3639, new_G3642, new_G3645,
    new_G3653, new_G3654, new_G3655, new_G3656, new_G763, new_G764,
    new_G803, new_G804, new_G1657, new_G1659, new_G2328, new_G2330,
    new_G1662, new_G2333, new_G657, new_G689;
  assign G144 = G141;
  assign G298 = G293;
  assign new_G4114 = G135 & G4115;
  assign new_G2825 = ~G2824;
  assign G973 = G3173;
  assign new_G3547 = ~G3546;
  assign new_G3549 = ~G3548;
  assign new_G3551 = ~G3550;
  assign new_G3553 = ~G3552;
  assign G594 = ~G545;
  assign G599 = ~G348;
  assign G600 = ~G366;
  assign G601 = G552 & G562;
  assign G602 = ~G549;
  assign G603 = ~G545;
  assign G604 = ~G545;
  assign G611 = ~G338;
  assign G612 = ~G358;
  assign new_G633 = ~G373 | ~G1;
  assign G810 = G141 & G145;
  assign new_G814 = ~G3173;
  assign new_G816 = ~new_G4114;
  assign new_G844 = new_G2825 & G27;
  assign new_G846 = G386 & G556;
  assign G848 = ~G245;
  assign G849 = ~G552;
  assign G850 = ~G562;
  assign G851 = ~G559;
  assign new_G852 = G552 & G556 & G386 & G559;
  assign new_G1502 = ~G1497;
  assign new_G1528 = G1689;
  assign new_G1552 = G1690;
  assign new_G1609 = G1689;
  assign new_G1633 = G1690;
  assign new_G1697 = G137;
  assign new_G1698 = G137;
  assign new_G1701 = G141;
  assign new_G2179 = ~G2174;
  assign new_G2203 = G1691;
  assign new_G2226 = G1694;
  assign new_G2281 = G1691;
  assign new_G2304 = G1694;
  assign new_G2361 = G254;
  assign new_G2370 = G251;
  assign new_G2382 = G251;
  assign new_G2393 = G248;
  assign new_G2405 = G248;
  assign new_G2418 = G4088;
  assign new_G2442 = G4087;
  assign new_G2476 = G4089;
  assign new_G2500 = G4090;
  assign new_G2533 = G210;
  assign new_G2537 = G210;
  assign new_G2541 = G218;
  assign new_G2545 = G218;
  assign new_G2549 = G226;
  assign new_G2553 = G226;
  assign new_G2557 = G234;
  assign new_G2561 = G234;
  assign new_G2627 = G257;
  assign new_G2631 = G257;
  assign new_G2635 = G265;
  assign new_G2639 = G265;
  assign new_G2643 = G273;
  assign new_G2647 = G273;
  assign new_G2651 = G281;
  assign new_G2655 = G281;
  assign new_G2721 = G335;
  assign new_G2734 = G335;
  assign new_G2816 = G206;
  assign new_G2822 = G27 & G31;
  assign new_G2826 = G1;
  assign new_G2828 = G2358;
  assign new_G2882 = G293;
  assign new_G2886 = G302;
  assign new_G2890 = G308;
  assign new_G2894 = G308;
  assign new_G2898 = G316;
  assign new_G2902 = G316;
  assign new_G2948 = G324;
  assign new_G2952 = G324;
  assign new_G2956 = G341;
  assign new_G2960 = G341;
  assign new_G2964 = G351;
  assign new_G2968 = G351;
  assign new_G3024 = G257;
  assign new_G3028 = G257;
  assign new_G3032 = G265;
  assign new_G3036 = G265;
  assign new_G3040 = G273;
  assign new_G3044 = G273;
  assign new_G3048 = G281;
  assign new_G3052 = G281;
  assign new_G3092 = G332;
  assign new_G3105 = G332;
  assign new_G3175 = G549;
  assign new_G3176 = G31 & G27;
  assign new_G3181 = ~G2358;
  assign new_G3204 = G324;
  assign new_G3208 = G324;
  assign new_G3212 = G341;
  assign new_G3216 = G341;
  assign new_G3220 = G351;
  assign new_G3224 = G351;
  assign new_G3256 = G293;
  assign new_G3260 = G302;
  assign new_G3264 = G308;
  assign new_G3268 = G308;
  assign new_G3272 = G316;
  assign new_G3276 = G316;
  assign new_G3302 = G361;
  assign new_G3314 = G361;
  assign new_G3354 = G210;
  assign new_G3358 = G210;
  assign new_G3362 = G218;
  assign new_G3366 = G218;
  assign new_G3370 = G226;
  assign new_G3374 = G226;
  assign new_G3378 = G234;
  assign new_G3382 = G234;
  assign new_G3440 = ~G324;
  assign new_G3554 = G242;
  assign new_G3555 = G242;
  assign new_G3556 = G254;
  assign new_G3558 = G4088;
  assign new_G3582 = G4087;
  assign new_G3616 = G4092;
  assign new_G3628 = G4091;
  assign new_G3660 = G4089;
  assign new_G3684 = G4090;
  assign new_G3721 = ~G3717;
  assign new_G3728 = ~G3724;
  assign new_G3737 = G4091;
  assign new_G3757 = G4092;
  assign new_G3795 = G4091;
  assign new_G3815 = G4092;
  assign new_G3972 = G4091;
  assign new_G3991 = G4092;
  assign new_G4030 = G4091;
  assign new_G4049 = G4092;
  assign new_G4110 = G299;
  assign new_G4119 = G446;
  assign new_G4127 = G457;
  assign new_G4135 = G468;
  assign new_G4143 = G422;
  assign new_G4151 = G435;
  assign new_G4159 = G389;
  assign new_G4167 = G400;
  assign new_G4175 = G411;
  assign new_G4183 = G374;
  assign new_G4188 = G4;
  assign new_G4276 = G446;
  assign new_G4284 = G457;
  assign new_G4292 = G468;
  assign new_G4300 = G435;
  assign new_G4308 = G389;
  assign new_G4316 = G400;
  assign new_G4324 = G411;
  assign new_G4332 = G422;
  assign new_G4340 = G374;
  assign new_G4631 = G479;
  assign new_G4639 = G490;
  assign new_G4647 = G503;
  assign new_G4655 = G514;
  assign new_G4663 = G523;
  assign new_G4671 = G534;
  assign new_G4676 = G54;
  assign new_G4764 = G479;
  assign new_G4772 = G503;
  assign new_G4780 = G514;
  assign new_G4788 = G523;
  assign new_G4796 = G534;
  assign new_G4804 = G490;
  assign new_G5082 = G361;
  assign new_G5085 = G369;
  assign new_G5090 = G341;
  assign new_G5093 = G351;
  assign new_G5098 = G308;
  assign new_G5101 = G316;
  assign new_G5108 = G293;
  assign new_G5111 = G302;
  assign new_G5332 = G281;
  assign new_G5335 = G289;
  assign new_G5340 = G265;
  assign new_G5343 = G273;
  assign new_G5348 = G234;
  assign new_G5351 = G257;
  assign new_G5356 = G218;
  assign new_G5359 = G226;
  assign new_G5369 = G210;
  assign G634 = ~new_G633;
  assign G815 = G136 & new_G814;
  assign G845 = ~new_G844;
  assign G847 = ~new_G846;
  assign G926 = new_G1697;
  assign G923 = new_G1701;
  assign G921 = new_G2826;
  assign new_G2979 = new_G3553 & G514;
  assign new_G2999 = new_G3547 | G514;
  assign G892 = new_G3175;
  assign G887 = new_G4110;
  assign G606 = ~new_G3175;
  assign new_G1580 = new_G1552 & G170 & new_G1528;
  assign new_G1586 = new_G1552 & G173 & new_G1528;
  assign new_G1592 = new_G1552 & G167 & new_G1528;
  assign new_G1598 = new_G1552 & G164 & new_G1528;
  assign new_G1604 = new_G1552 & G161 & new_G1528;
  assign G656 = ~new_G2822 | ~G140;
  assign new_G1668 = new_G1633 & G185 & new_G1609;
  assign new_G1674 = new_G1633 & G158 & new_G1609;
  assign new_G1680 = new_G1633 & G152 & new_G1609;
  assign new_G1686 = new_G1633 & G146 & new_G1609;
  assign new_G2254 = new_G2226 & G170 & new_G2203;
  assign new_G2260 = new_G2226 & G173 & new_G2203;
  assign new_G2266 = new_G2226 & G167 & new_G2203;
  assign new_G2272 = new_G2226 & G164 & new_G2203;
  assign new_G2278 = new_G2226 & G161 & new_G2203;
  assign new_G2339 = new_G2304 & G185 & new_G2281;
  assign new_G2345 = new_G2304 & G158 & new_G2281;
  assign new_G2351 = new_G2304 & G152 & new_G2281;
  assign new_G2357 = new_G2304 & G146 & new_G2281;
  assign new_G711 = new_G3684 & G106 & new_G3660;
  assign new_G721 = new_G2442 & G61 & new_G2418;
  assign new_G726 = new_G3582 & G106 & new_G3558;
  assign new_G731 = new_G3582 & G49 & new_G3558;
  assign new_G736 = new_G3582 & G103 & new_G3558;
  assign new_G741 = new_G3582 & G40 & new_G3558;
  assign new_G746 = new_G3582 & G37 & new_G3558;
  assign new_G751 = new_G2442 & G20 & new_G2418;
  assign new_G756 = new_G2442 & G17 & new_G2418;
  assign new_G761 = new_G2442 & G70 & new_G2418;
  assign new_G766 = new_G2442 & G64 & new_G2418;
  assign new_G771 = new_G3684 & G49 & new_G3660;
  assign new_G776 = new_G3684 & G103 & new_G3660;
  assign new_G781 = new_G3684 & G40 & new_G3660;
  assign new_G786 = new_G3684 & G37 & new_G3660;
  assign new_G791 = new_G2500 & G20 & new_G2476;
  assign new_G796 = new_G2500 & G17 & new_G2476;
  assign new_G801 = new_G2500 & G70 & new_G2476;
  assign new_G806 = new_G2500 & G64 & new_G2476;
  assign G809 = ~new_G2822;
  assign new_G3734 = G3717 & G123 & new_G3728;
  assign new_G842 = new_G3795 & new_G3815;
  assign new_G858 = new_G2500 & G61 & new_G2476;
  assign new_G881 = new_G3737 & new_G3757;
  assign new_G4123 = ~new_G4119;
  assign new_G4131 = ~new_G4127;
  assign new_G4139 = ~new_G4135;
  assign new_G4147 = ~new_G4143;
  assign new_G4155 = ~new_G4151;
  assign new_G4163 = ~new_G4159;
  assign new_G4171 = ~new_G4167;
  assign new_G4179 = ~new_G4175;
  assign new_G4187 = ~new_G4183;
  assign new_G4194 = ~new_G4188;
  assign new_G4282 = ~new_G4276;
  assign new_G4290 = ~new_G4284;
  assign new_G4298 = ~new_G4292;
  assign new_G4306 = ~new_G4300;
  assign new_G4314 = ~new_G4308;
  assign new_G4322 = ~new_G4316;
  assign new_G4330 = ~new_G4324;
  assign new_G4338 = ~new_G4332;
  assign new_G4346 = ~new_G4340;
  assign new_G1526 = new_G1697;
  assign new_G1540 = ~new_G1528;
  assign new_G1564 = ~new_G1552;
  assign new_G1606 = new_G1697;
  assign new_G1621 = ~new_G1609;
  assign new_G1645 = ~new_G1633;
  assign new_G1661 = new_G1633 & G179 & new_G1609;
  assign new_G1688 = new_G2826;
  assign new_G4635 = ~new_G4631;
  assign new_G4643 = ~new_G4639;
  assign new_G4651 = ~new_G4647;
  assign new_G4659 = ~new_G4655;
  assign new_G4667 = ~new_G4663;
  assign new_G4675 = ~new_G4671;
  assign new_G4682 = ~new_G4676;
  assign new_G4770 = ~new_G4764;
  assign new_G4778 = ~new_G4772;
  assign new_G4786 = ~new_G4780;
  assign new_G4794 = ~new_G4788;
  assign new_G4802 = ~new_G4796;
  assign new_G4810 = ~new_G4804;
  assign new_G2202 = new_G1698;
  assign new_G2215 = ~new_G2203;
  assign new_G2238 = ~new_G2226;
  assign new_G2279 = new_G1698;
  assign new_G2293 = ~new_G2281;
  assign new_G2316 = ~new_G2304;
  assign new_G2332 = new_G2304 & G179 & new_G2281;
  assign new_G2430 = ~new_G2418;
  assign new_G2454 = ~new_G2442;
  assign new_G2488 = ~new_G2476;
  assign new_G2512 = ~new_G2500;
  assign new_G2536 = ~new_G2533;
  assign new_G2540 = ~new_G2537;
  assign new_G2544 = ~new_G2541;
  assign new_G2548 = ~new_G2545;
  assign new_G2552 = ~new_G2549;
  assign new_G2556 = ~new_G2553;
  assign new_G2560 = ~new_G2557;
  assign new_G2564 = ~new_G2561;
  assign new_G2566 = new_G2537 & new_G3553 & G457;
  assign new_G2572 = new_G2545 & new_G3553 & G468;
  assign new_G2578 = new_G2553 & new_G3553 & G422;
  assign new_G2584 = new_G2561 & new_G3553 & G435;
  assign new_G2590 = new_G3547 & new_G2533;
  assign new_G2595 = new_G3547 & new_G2541;
  assign new_G2600 = new_G3547 & new_G2549;
  assign new_G2605 = new_G3547 & new_G2557;
  assign new_G2630 = ~new_G2627;
  assign new_G2634 = ~new_G2631;
  assign new_G2638 = ~new_G2635;
  assign new_G2642 = ~new_G2639;
  assign new_G2646 = ~new_G2643;
  assign new_G2650 = ~new_G2647;
  assign new_G2654 = ~new_G2651;
  assign new_G2658 = ~new_G2655;
  assign new_G2660 = new_G2631 & new_G3553 & G389;
  assign new_G2666 = new_G2639 & new_G3553 & G400;
  assign new_G2672 = new_G2647 & new_G3553 & G411;
  assign new_G2678 = new_G2655 & new_G3553 & G374;
  assign new_G2684 = new_G3547 & new_G2627;
  assign new_G2689 = new_G3547 & new_G2635;
  assign new_G2694 = new_G3547 & new_G2643;
  assign new_G2699 = new_G3547 & new_G2651;
  assign new_G2728 = ~new_G2721;
  assign new_G2741 = ~new_G2734;
  assign new_G2748 = G292 & new_G2721;
  assign new_G2750 = G288 & new_G2721;
  assign new_G2752 = G280 & new_G2721;
  assign new_G2754 = G272 & new_G2721;
  assign new_G2756 = G264 & new_G2721;
  assign new_G2758 = G241 & new_G2734;
  assign new_G2760 = G233 & new_G2734;
  assign new_G2762 = G225 & new_G2734;
  assign new_G2764 = G217 & new_G2734;
  assign new_G2766 = G209 & new_G2734;
  assign new_G2827 = new_G1701;
  assign new_G2838 = ~new_G2828;
  assign new_G2847 = ~new_G2822;
  assign new_G2885 = ~new_G2882;
  assign new_G2889 = ~new_G2886;
  assign new_G2893 = ~new_G2890;
  assign new_G2897 = ~new_G2894;
  assign new_G2901 = ~new_G2898;
  assign new_G2905 = ~new_G2902;
  assign new_G2906 = new_G2393 & new_G2886;
  assign new_G2909 = new_G2894 & new_G2393 & G479;
  assign new_G2913 = new_G2902 & new_G2393 & G490;
  assign new_G2918 = new_G3554 & new_G2882;
  assign new_G2922 = new_G3554 & new_G2890;
  assign new_G2927 = new_G3554 & new_G2898;
  assign new_G2951 = ~new_G2948;
  assign new_G2955 = ~new_G2952;
  assign new_G2959 = ~new_G2956;
  assign new_G2963 = ~new_G2960;
  assign new_G2967 = ~new_G2964;
  assign new_G2971 = ~new_G2968;
  assign new_G2973 = new_G2952 & new_G3553 & G503;
  assign new_G2980 = ~new_G2979;
  assign new_G2982 = new_G2960 & new_G3553 & G523;
  assign new_G2988 = new_G2968 & new_G3553 & G534;
  assign new_G2994 = new_G3547 & new_G2948;
  assign new_G3001 = new_G3547 & new_G2956;
  assign new_G3006 = new_G3547 & new_G2964;
  assign new_G3027 = ~new_G3024;
  assign new_G3031 = ~new_G3028;
  assign new_G3035 = ~new_G3032;
  assign new_G3039 = ~new_G3036;
  assign new_G3043 = ~new_G3040;
  assign new_G3047 = ~new_G3044;
  assign new_G3051 = ~new_G3048;
  assign new_G3055 = ~new_G3052;
  assign new_G3056 = new_G3028 & new_G2393 & G389;
  assign new_G3060 = new_G3036 & new_G2393 & G400;
  assign new_G3064 = new_G3044 & new_G2393 & G411;
  assign new_G3068 = new_G3052 & new_G2393 & G374;
  assign new_G3073 = new_G3554 & new_G3024;
  assign new_G3078 = new_G3554 & new_G3032;
  assign new_G3083 = new_G3554 & new_G3040;
  assign new_G3088 = new_G3554 & new_G3048;
  assign new_G3099 = ~new_G3092;
  assign new_G3112 = ~new_G3105;
  assign new_G3119 = G372 & new_G3092;
  assign new_G3121 = G366 & new_G3092;
  assign new_G3123 = G358 & new_G3092;
  assign new_G3125 = G348 & new_G3092;
  assign new_G3126 = G338 & new_G3092;
  assign new_G3128 = G331 & new_G3105;
  assign new_G3130 = G323 & new_G3105;
  assign new_G3132 = G315 & new_G3105;
  assign new_G3134 = G307 & new_G3105;
  assign new_G3136 = G299 & new_G3105;
  assign new_G3187 = ~new_G3181;
  assign new_G3193 = G83 & new_G3181;
  assign new_G3196 = G86 & new_G3181;
  assign new_G3199 = G88 & new_G3181;
  assign new_G3202 = G88 & new_G3181;
  assign new_G3207 = ~new_G3204;
  assign new_G3211 = ~new_G3208;
  assign new_G3215 = ~new_G3212;
  assign new_G3219 = ~new_G3216;
  assign new_G3223 = ~new_G3220;
  assign new_G3227 = ~new_G3224;
  assign new_G3228 = new_G3208 & new_G2405 & G503;
  assign new_G3232 = new_G2405 & G514;
  assign new_G3234 = new_G3216 & new_G2405 & G523;
  assign new_G3238 = new_G3224 & new_G2405 & G534;
  assign new_G3243 = new_G3555 & new_G3204;
  assign new_G3247 = new_G3555 | G514;
  assign new_G3249 = new_G3555 & new_G3212;
  assign new_G3253 = new_G3555 & new_G3220;
  assign new_G3259 = ~new_G3256;
  assign new_G3263 = ~new_G3260;
  assign new_G3267 = ~new_G3264;
  assign new_G3271 = ~new_G3268;
  assign new_G3275 = ~new_G3272;
  assign new_G3279 = ~new_G3276;
  assign new_G3280 = new_G2405 & new_G3260;
  assign new_G3283 = new_G3268 & new_G2405 & G479;
  assign new_G3287 = new_G3276 & new_G2405 & G490;
  assign new_G3292 = new_G3555 & new_G3256;
  assign new_G3295 = new_G3555 & new_G3264;
  assign new_G3299 = new_G3555 & new_G3272;
  assign new_G3305 = ~new_G3302;
  assign new_G3306 = new_G2816;
  assign new_G3310 = new_G2816;
  assign new_G3317 = ~new_G3314;
  assign new_G3318 = new_G2816;
  assign new_G3322 = new_G2816;
  assign new_G3326 = new_G2405 & new_G3302;
  assign new_G3333 = new_G2405 & new_G3314;
  assign new_G3357 = ~new_G3354;
  assign new_G3361 = ~new_G3358;
  assign new_G3365 = ~new_G3362;
  assign new_G3369 = ~new_G3366;
  assign new_G3373 = ~new_G3370;
  assign new_G3377 = ~new_G3374;
  assign new_G3381 = ~new_G3378;
  assign new_G3385 = ~new_G3382;
  assign new_G3386 = new_G3358 & new_G2393 & G457;
  assign new_G3390 = new_G3366 & new_G2393 & G468;
  assign new_G3394 = new_G3374 & new_G2393 & G422;
  assign new_G3398 = new_G3382 & new_G2393 & G435;
  assign new_G3403 = new_G3554 & new_G3354;
  assign new_G3408 = new_G3554 & new_G3362;
  assign new_G3413 = new_G3554 & new_G3370;
  assign new_G3418 = new_G3554 & new_G3378;
  assign new_G5088 = ~new_G5082;
  assign new_G5089 = ~new_G5085;
  assign new_G5096 = ~new_G5090;
  assign new_G5097 = ~new_G5093;
  assign new_G3489 = new_G3440;
  assign new_G3493 = new_G3440;
  assign new_G3570 = ~new_G3558;
  assign new_G3594 = ~new_G3582;
  assign new_G3622 = ~new_G3616;
  assign new_G3632 = ~new_G3628;
  assign new_G3637 = G97 & new_G3616;
  assign new_G3640 = G94 & new_G3616;
  assign new_G3643 = G97 & new_G3616;
  assign new_G3646 = G94 & new_G3616;
  assign new_G3672 = ~new_G3660;
  assign new_G3696 = ~new_G3684;
  assign new_G3745 = ~new_G3737;
  assign new_G3765 = ~new_G3757;
  assign new_G3803 = ~new_G3795;
  assign new_G3823 = ~new_G3815;
  assign new_G5338 = ~new_G5332;
  assign new_G5339 = ~new_G5335;
  assign new_G5346 = ~new_G5340;
  assign new_G5347 = ~new_G5343;
  assign new_G5354 = ~new_G5348;
  assign new_G5355 = ~new_G5351;
  assign new_G3979 = ~new_G3972;
  assign new_G3998 = ~new_G3991;
  assign new_G4037 = ~new_G4030;
  assign new_G4056 = ~new_G4049;
  assign new_G4094 = new_G4110;
  assign new_G5104 = ~new_G5098;
  assign new_G5105 = ~new_G5101;
  assign new_G5114 = ~new_G5108;
  assign new_G5115 = ~new_G5111;
  assign new_G5362 = ~new_G5356;
  assign new_G5363 = ~new_G5359;
  assign new_G5366 = new_G2816;
  assign new_G5373 = ~new_G5369;
  assign G993 = new_G1688;
  assign G978 = new_G1688;
  assign G949 = new_G1688;
  assign G939 = new_G1688;
  assign new_G2568 = new_G2540 & G457 & new_G3551;
  assign new_G2574 = new_G2548 & G468 & new_G3551;
  assign new_G2580 = new_G2556 & G422 & new_G3551;
  assign new_G2586 = new_G2564 & G435 & new_G3551;
  assign new_G2592 = new_G3549 & new_G2536;
  assign new_G2597 = new_G3549 & new_G2544;
  assign new_G2602 = new_G3549 & new_G2552;
  assign new_G2607 = new_G3549 & new_G2560;
  assign new_G2662 = new_G2634 & G389 & new_G3551;
  assign new_G2668 = new_G2642 & G400 & new_G3551;
  assign new_G2674 = new_G2650 & G411 & new_G3551;
  assign new_G2680 = new_G2658 & G374 & new_G3551;
  assign new_G2686 = new_G3549 & new_G2630;
  assign new_G2691 = new_G3549 & new_G2638;
  assign new_G2696 = new_G3549 & new_G2646;
  assign new_G2701 = new_G3549 & new_G2654;
  assign new_G2907 = new_G2370 & new_G2889;
  assign new_G2910 = new_G2897 & G479 & new_G2370;
  assign new_G2914 = new_G2905 & G490 & new_G2370;
  assign new_G2920 = new_G3556 & new_G2885;
  assign new_G2924 = new_G3556 & new_G2893;
  assign new_G2929 = new_G3556 & new_G2901;
  assign new_G2975 = new_G2955 & G503 & new_G3551;
  assign new_G2984 = new_G2963 & G523 & new_G3551;
  assign new_G2990 = new_G2971 & G534 & new_G3551;
  assign new_G2996 = new_G3549 & new_G2951;
  assign new_G3003 = new_G3549 & new_G2959;
  assign new_G3008 = new_G3549 & new_G2967;
  assign new_G3015 = new_G2980 & new_G2999;
  assign new_G3057 = new_G3031 & G389 & new_G2370;
  assign new_G3061 = new_G3039 & G400 & new_G2370;
  assign new_G3065 = new_G3047 & G411 & new_G2370;
  assign new_G3069 = new_G3055 & G374 & new_G2370;
  assign new_G3075 = new_G3556 & new_G3027;
  assign new_G3080 = new_G3556 & new_G3035;
  assign new_G3085 = new_G3556 & new_G3043;
  assign new_G3090 = new_G3556 & new_G3051;
  assign new_G3229 = new_G3211 & G503 & new_G2382;
  assign new_G3233 = ~new_G3232;
  assign new_G3235 = new_G3219 & G523 & new_G2382;
  assign new_G3239 = new_G3227 & G534 & new_G2382;
  assign new_G3244 = new_G2361 & new_G3207;
  assign new_G3250 = new_G2361 & new_G3215;
  assign new_G3254 = new_G2361 & new_G3223;
  assign new_G3281 = new_G2382 & new_G3263;
  assign new_G3284 = new_G3271 & G479 & new_G2382;
  assign new_G3288 = new_G3279 & G490 & new_G2382;
  assign new_G3293 = new_G2361 & new_G3259;
  assign new_G3296 = new_G2361 & new_G3267;
  assign new_G3300 = new_G2361 & new_G3275;
  assign new_G3327 = new_G2382 & new_G3305;
  assign new_G3334 = new_G2382 & new_G3317;
  assign new_G3387 = new_G3361 & G457 & new_G2370;
  assign new_G3391 = new_G3369 & G468 & new_G2370;
  assign new_G3395 = new_G3377 & G422 & new_G2370;
  assign new_G3399 = new_G3385 & G435 & new_G2370;
  assign new_G3405 = new_G3556 & new_G3357;
  assign new_G3410 = new_G3556 & new_G3365;
  assign new_G3415 = new_G3556 & new_G3373;
  assign new_G3420 = new_G3556 & new_G3381;
  assign new_G3422 = ~new_G5085 | ~new_G5088;
  assign new_G3423 = ~new_G5082 | ~new_G5089;
  assign new_G3431 = ~new_G5093 | ~new_G5096;
  assign new_G3432 = ~new_G5090 | ~new_G5097;
  assign new_G3895 = ~new_G5335 | ~new_G5338;
  assign new_G3896 = ~new_G5332 | ~new_G5339;
  assign new_G3904 = ~new_G5343 | ~new_G5346;
  assign new_G3905 = ~new_G5340 | ~new_G5347;
  assign new_G3913 = ~new_G5351 | ~new_G5354;
  assign new_G3914 = ~new_G5348 | ~new_G5355;
  assign G889 = new_G4094;
  assign new_G5106 = ~new_G5101 | ~new_G5104;
  assign new_G5107 = ~new_G5098 | ~new_G5105;
  assign new_G5116 = ~new_G5111 | ~new_G5114;
  assign new_G5117 = ~new_G5108 | ~new_G5115;
  assign new_G5364 = ~new_G5359 | ~new_G5362;
  assign new_G5365 = ~new_G5356 | ~new_G5363;
  assign G593 = ~new_G4094;
  assign new_G2880 = new_G2838 & new_G2847;
  assign new_G2881 = new_G2828 & new_G2847;
  assign new_G1579 = new_G1552 & G200 & new_G1540;
  assign new_G1585 = new_G1552 & G203 & new_G1540;
  assign new_G1591 = new_G1552 & G197 & new_G1540;
  assign new_G1597 = new_G1552 & G194 & new_G1540;
  assign new_G1603 = new_G1552 & G191 & new_G1540;
  assign new_G1667 = new_G1633 & G182 & new_G1621;
  assign new_G1673 = new_G1633 & G188 & new_G1621;
  assign new_G1679 = new_G1633 & G155 & new_G1621;
  assign new_G1685 = new_G1633 & G149 & new_G1621;
  assign new_G2876 = new_G2838 & new_G2847;
  assign new_G2877 = new_G2828 & new_G2847;
  assign new_G2253 = new_G2226 & G200 & new_G2215;
  assign new_G2259 = new_G2226 & G203 & new_G2215;
  assign new_G2265 = new_G2226 & G197 & new_G2215;
  assign new_G2271 = new_G2226 & G194 & new_G2215;
  assign new_G2277 = new_G2226 & G191 & new_G2215;
  assign new_G2338 = new_G2304 & G182 & new_G2293;
  assign new_G2344 = new_G2304 & G188 & new_G2293;
  assign new_G2350 = new_G2304 & G155 & new_G2293;
  assign new_G2356 = new_G2304 & G149 & new_G2293;
  assign new_G2868 = new_G2838 & new_G2847;
  assign new_G2869 = new_G2828 & new_G2847;
  assign new_G710 = new_G3684 & G109 & new_G3672;
  assign new_G2872 = new_G2838 & new_G2847;
  assign new_G2873 = new_G2828 & new_G2847;
  assign new_G720 = new_G2442 & G11 & new_G2430;
  assign new_G725 = new_G3582 & G109 & new_G3570;
  assign new_G730 = new_G3582 & G46 & new_G3570;
  assign new_G735 = new_G3582 & G100 & new_G3570;
  assign new_G740 = new_G3582 & G91 & new_G3570;
  assign new_G745 = new_G3582 & G43 & new_G3570;
  assign new_G750 = new_G2442 & G76 & new_G2430;
  assign new_G755 = new_G2442 & G73 & new_G2430;
  assign new_G760 = new_G2442 & G67 & new_G2430;
  assign new_G765 = new_G2442 & G14 & new_G2430;
  assign new_G770 = new_G3684 & G46 & new_G3672;
  assign new_G775 = new_G3684 & G100 & new_G3672;
  assign new_G780 = new_G3684 & G91 & new_G3672;
  assign new_G785 = new_G3684 & G43 & new_G3672;
  assign new_G790 = new_G2500 & G76 & new_G2488;
  assign new_G795 = new_G2500 & G73 & new_G2488;
  assign new_G800 = new_G2500 & G67 & new_G2488;
  assign new_G805 = new_G2500 & G14 & new_G2488;
  assign new_G841 = new_G3815 & G120 & new_G3803;
  assign new_G857 = new_G2500 & G11 & new_G2488;
  assign new_G880 = new_G3757 & G118 & new_G3745;
  assign new_G1660 = new_G1633 & G176 & new_G1621;
  assign new_G2331 = new_G2304 & G176 & new_G2293;
  assign new_G2569 = new_G2566 | new_G2568;
  assign new_G2575 = new_G2572 | new_G2574;
  assign new_G2581 = new_G2578 | new_G2580;
  assign new_G2587 = new_G2584 | new_G2586;
  assign new_G2593 = G457 | new_G2590 | new_G2592;
  assign new_G2598 = G468 | new_G2595 | new_G2597;
  assign new_G2603 = G422 | new_G2600 | new_G2602;
  assign new_G2608 = G435 | new_G2605 | new_G2607;
  assign new_G2663 = new_G2660 | new_G2662;
  assign new_G2669 = new_G2666 | new_G2668;
  assign new_G2675 = new_G2672 | new_G2674;
  assign new_G2681 = new_G2678 | new_G2680;
  assign new_G2687 = G389 | new_G2684 | new_G2686;
  assign new_G2692 = G400 | new_G2689 | new_G2691;
  assign new_G2697 = G411 | new_G2694 | new_G2696;
  assign new_G2702 = G374 | new_G2699 | new_G2701;
  assign new_G2747 = G289 & new_G2728;
  assign new_G2749 = G281 & new_G2728;
  assign new_G2751 = G273 & new_G2728;
  assign new_G2753 = G265 & new_G2728;
  assign new_G2755 = G257 & new_G2728;
  assign new_G2757 = G234 & new_G2741;
  assign new_G2759 = G226 & new_G2741;
  assign new_G2761 = G218 & new_G2741;
  assign new_G2763 = G210 & new_G2741;
  assign new_G2765 = G206 & new_G2741;
  assign new_G2857 = ~new_G2847;
  assign new_G2908 = new_G2906 | new_G2907;
  assign new_G2911 = new_G2909 | new_G2910;
  assign new_G2915 = new_G2913 | new_G2914;
  assign new_G2925 = G479 | new_G2922 | new_G2924;
  assign new_G2930 = G490 | new_G2927 | new_G2929;
  assign new_G2933 = new_G2918 | new_G2920;
  assign new_G2976 = new_G2973 | new_G2975;
  assign new_G2985 = new_G2982 | new_G2984;
  assign new_G2991 = new_G2988 | new_G2990;
  assign new_G2997 = G503 | new_G2994 | new_G2996;
  assign new_G3004 = G523 | new_G3001 | new_G3003;
  assign new_G3009 = G534 | new_G3006 | new_G3008;
  assign new_G3058 = new_G3056 | new_G3057;
  assign new_G3062 = new_G3060 | new_G3061;
  assign new_G3066 = new_G3064 | new_G3065;
  assign new_G3070 = new_G3068 | new_G3069;
  assign new_G3076 = G389 | new_G3073 | new_G3075;
  assign new_G3081 = G400 | new_G3078 | new_G3080;
  assign new_G3086 = G411 | new_G3083 | new_G3085;
  assign new_G3091 = G374 | new_G3088 | new_G3090;
  assign new_G3118 = G369 & new_G3099;
  assign new_G3120 = G361 & new_G3099;
  assign new_G3122 = G351 & new_G3099;
  assign new_G3124 = G341 & new_G3099;
  assign new_G3127 = G324 & new_G3112;
  assign new_G3129 = G316 & new_G3112;
  assign new_G3131 = G308 & new_G3112;
  assign new_G3133 = G302 & new_G3112;
  assign new_G3135 = G293 & new_G3112;
  assign new_G3147 = new_G3099 | new_G3126;
  assign new_G3192 = G83 & new_G3187;
  assign new_G3195 = G87 & new_G3187;
  assign new_G3198 = G34 & new_G3187;
  assign new_G3201 = G34 & new_G3187;
  assign new_G3230 = new_G3228 | new_G3229;
  assign new_G3236 = new_G3234 | new_G3235;
  assign new_G3240 = new_G3238 | new_G3239;
  assign new_G3245 = G503 | new_G3243 | new_G3244;
  assign new_G3251 = G523 | new_G3249 | new_G3250;
  assign new_G3255 = G534 | new_G3253 | new_G3254;
  assign new_G3282 = new_G3280 | new_G3281;
  assign new_G3285 = new_G3283 | new_G3284;
  assign new_G3289 = new_G3287 | new_G3288;
  assign new_G3297 = G479 | new_G3295 | new_G3296;
  assign new_G3301 = G490 | new_G3299 | new_G3300;
  assign new_G3309 = ~new_G3306;
  assign new_G3313 = ~new_G3310;
  assign new_G3321 = ~new_G3318;
  assign new_G3325 = ~new_G3322;
  assign new_G3328 = new_G3326 | new_G3327;
  assign new_G3329 = new_G3310 & new_G2405 & G446;
  assign new_G3335 = new_G3333 | new_G3334;
  assign new_G3336 = new_G3322 & new_G2405 & G446;
  assign new_G3341 = new_G3555 & new_G3306;
  assign new_G3345 = new_G3555 & new_G3318;
  assign new_G3388 = new_G3386 | new_G3387;
  assign new_G3392 = new_G3390 | new_G3391;
  assign new_G3396 = new_G3394 | new_G3395;
  assign new_G3400 = new_G3398 | new_G3399;
  assign new_G3406 = G457 | new_G3403 | new_G3405;
  assign new_G3411 = G468 | new_G3408 | new_G3410;
  assign new_G3416 = G422 | new_G3413 | new_G3415;
  assign new_G3421 = G435 | new_G3418 | new_G3420;
  assign new_G3424 = ~new_G3422 | ~new_G3423;
  assign new_G3433 = ~new_G3431 | ~new_G3432;
  assign new_G3492 = ~new_G3489;
  assign new_G3496 = ~new_G3493;
  assign new_G3780 = new_G3757 & G117 & new_G3745;
  assign new_G3783 = new_G3757 & G126 & new_G3745;
  assign new_G3786 = new_G3757 & G127 & new_G3745;
  assign new_G3789 = new_G3757 & G128 & new_G3745;
  assign new_G3838 = new_G3815 & G131 & new_G3803;
  assign new_G3841 = new_G3815 & G129 & new_G3803;
  assign new_G3844 = new_G3815 & G119 & new_G3803;
  assign new_G3847 = new_G3815 & G130 & new_G3803;
  assign new_G3897 = ~new_G3895 | ~new_G3896;
  assign new_G3906 = ~new_G3904 | ~new_G3905;
  assign new_G3915 = ~new_G3913 | ~new_G3914;
  assign new_G4011 = new_G3991 & G122 & new_G3979;
  assign new_G4014 = new_G3991 & G113 & new_G3979;
  assign new_G4017 = new_G3991 & G53 & new_G3979;
  assign new_G4020 = new_G3991 & G114 & new_G3979;
  assign new_G4023 = new_G3991 & G115 & new_G3979;
  assign new_G4069 = new_G4049 & G52 & new_G4037;
  assign new_G4072 = new_G4049 & G112 & new_G4037;
  assign new_G4075 = new_G4049 & G116 & new_G4037;
  assign new_G4078 = new_G4049 & G121 & new_G4037;
  assign new_G4081 = new_G4049 & G123 & new_G4037;
  assign new_G5206 = ~new_G5116 | ~new_G5117;
  assign new_G5209 = ~new_G5106 | ~new_G5107;
  assign new_G5307 = new_G3233 & new_G3247;
  assign new_G5322 = new_G3292 | new_G3293;
  assign new_G5372 = ~new_G5366;
  assign new_G5375 = ~new_G5366 | ~new_G5373;
  assign new_G5399 = ~new_G5364 | ~new_G5365;
  assign new_G2813 = ~new_G3015;
  assign new_G3197 = new_G3195 | new_G3196;
  assign new_G3200 = new_G3198 | new_G3199;
  assign new_G3203 = new_G3201 | new_G3202;
  assign new_G3194 = new_G3192 | new_G3193;
  assign new_G2570 = ~new_G2569;
  assign new_G2576 = ~new_G2575;
  assign new_G2582 = ~new_G2581;
  assign new_G2588 = ~new_G2587;
  assign new_G2664 = ~new_G2663;
  assign new_G2670 = ~new_G2669;
  assign new_G2676 = ~new_G2675;
  assign new_G2682 = ~new_G2681;
  assign new_G2767 = new_G2749 | new_G2750;
  assign new_G2772 = new_G2751 | new_G2752;
  assign new_G2776 = new_G2753 | new_G2754;
  assign new_G2780 = new_G2755 | new_G2756;
  assign new_G2784 = new_G2757 | new_G2758;
  assign new_G2788 = new_G2759 | new_G2760;
  assign new_G2794 = new_G2761 | new_G2762;
  assign new_G2798 = new_G2763 | new_G2764;
  assign new_G2802 = new_G2765 | new_G2766;
  assign new_G2912 = ~new_G2911;
  assign new_G2916 = ~new_G2915;
  assign new_G2936 = ~new_G2908;
  assign new_G2977 = ~new_G2976;
  assign new_G2986 = ~new_G2985;
  assign new_G2992 = ~new_G2991;
  assign new_G3059 = ~new_G3058;
  assign new_G3063 = ~new_G3062;
  assign new_G3067 = ~new_G3066;
  assign new_G3071 = ~new_G3070;
  assign new_G3137 = new_G3120 | new_G3121;
  assign new_G3139 = new_G3122 | new_G3123;
  assign new_G3143 = new_G3124 | new_G3125;
  assign new_G3151 = new_G3127 | new_G3128;
  assign new_G3155 = new_G3129 | new_G3130;
  assign new_G3161 = new_G3131 | new_G3132;
  assign new_G3165 = new_G3133 | new_G3134;
  assign new_G3167 = new_G3135 | new_G3136;
  assign new_G3231 = ~new_G3230;
  assign new_G3237 = ~new_G3236;
  assign new_G3241 = ~new_G3240;
  assign new_G3286 = ~new_G3285;
  assign new_G3290 = ~new_G3289;
  assign new_G3330 = new_G3313 & G446 & new_G2382;
  assign new_G3337 = new_G3325 & G446 & new_G2382;
  assign new_G3342 = new_G2361 & new_G3309;
  assign new_G3346 = new_G2361 & new_G3321;
  assign new_G3348 = ~new_G3328;
  assign new_G3352 = ~new_G3335;
  assign new_G3389 = ~new_G3388;
  assign new_G3393 = ~new_G3392;
  assign new_G3397 = ~new_G3396;
  assign new_G3401 = ~new_G3400;
  assign new_G3845 = new_G3823 & new_G3015 & new_G3803;
  assign new_G5126 = new_G3118 | new_G3119;
  assign new_G5178 = new_G2747 | new_G2748;
  assign new_G5325 = ~new_G3282;
  assign new_G5374 = ~new_G5369 | ~new_G5372;
  assign new_G2810 = ~new_G2933;
  assign new_G635 = new_G3197 & new_G3176;
  assign new_G2878 = new_G2857 & G24 & new_G2838;
  assign new_G2879 = new_G2857 & G25 & new_G2828;
  assign new_G2874 = new_G2857 & G26 & new_G2838;
  assign new_G2875 = new_G2857 & G81 & new_G2828;
  assign new_G703 = new_G3200 & new_G3176;
  assign new_G2866 = new_G2857 & G79 & new_G2838;
  assign new_G2867 = new_G2857 & G23 & new_G2828;
  assign new_G2870 = new_G2857 & G82 & new_G2838;
  assign new_G2871 = new_G2857 & G80 & new_G2828;
  assign new_G716 = new_G3203 & new_G3176;
  assign new_G819 = new_G3194 & new_G3176;
  assign new_G1789 = new_G3147 & G514;
  assign new_G2036 = G514 & new_G3147;
  assign new_G2611 = new_G2570 & new_G2593;
  assign new_G2615 = new_G2576 & new_G2598;
  assign new_G2619 = new_G2582 & new_G2603;
  assign new_G2623 = new_G2588 & new_G2608;
  assign new_G2705 = new_G2664 & new_G2687;
  assign new_G2709 = new_G2670 & new_G2692;
  assign new_G2713 = new_G2676 & new_G2697;
  assign new_G2717 = new_G2682 & new_G2702;
  assign new_G2939 = new_G2912 & new_G2925;
  assign new_G2942 = new_G2916 & new_G2930;
  assign new_G2945 = new_G2933;
  assign new_G3012 = new_G2977 & new_G2997;
  assign new_G3018 = new_G2986 & new_G3004;
  assign new_G3021 = new_G2992 & new_G3009;
  assign new_G3331 = new_G3329 | new_G3330;
  assign new_G3338 = new_G3336 | new_G3337;
  assign new_G3343 = G446 | new_G3341 | new_G3342;
  assign new_G3347 = G446 | new_G3345 | new_G3346;
  assign new_G3428 = ~new_G3424;
  assign new_G3437 = ~new_G3433;
  assign new_G3514 = new_G3489 & new_G3433 & new_G3424;
  assign new_G3836 = new_G3823 & new_G3352 & new_G3803;
  assign new_G3852 = new_G3071 & new_G3091;
  assign new_G5311 = ~new_G5307;
  assign new_G3901 = ~new_G3897;
  assign new_G3910 = ~new_G3906;
  assign new_G3934 = new_G3915;
  assign new_G3938 = new_G3915;
  assign new_G4652 = new_G3147;
  assign new_G4783 = new_G3147;
  assign new_G5137 = new_G3147;
  assign new_G5212 = ~new_G5206;
  assign new_G5213 = ~new_G5209;
  assign new_G5260 = new_G3063 & new_G3081;
  assign new_G5263 = new_G3067 & new_G3086;
  assign new_G5268 = new_G3401 & new_G3421;
  assign new_G5271 = new_G3059 & new_G3076;
  assign new_G5276 = new_G3393 & new_G3411;
  assign new_G5279 = new_G3397 & new_G3416;
  assign new_G5289 = new_G3389 & new_G3406;
  assign new_G5296 = new_G3237 & new_G3251;
  assign new_G5299 = new_G3241 & new_G3255;
  assign new_G5304 = new_G3231 & new_G3245;
  assign new_G5312 = new_G3286 & new_G3297;
  assign new_G5315 = new_G3290 & new_G3301;
  assign new_G5328 = ~new_G5322;
  assign new_G5396 = ~new_G5374 | ~new_G5375;
  assign new_G5403 = ~new_G5399;
  assign new_G1286 = G446 & new_G2802;
  assign new_G2809 = ~new_G2936;
  assign new_G597 = ~new_G3348;
  assign new_G1031 = new_G2802 & G446;
  assign G636 = ~new_G635;
  assign new_G637 = new_G2881 | new_G2880 | new_G2878 | new_G2879;
  assign new_G671 = new_G2877 | new_G2876 | new_G2874 | new_G2875;
  assign G704 = ~new_G703;
  assign new_G705 = new_G2869 | new_G2868 | new_G2866 | new_G2867;
  assign new_G713 = new_G2873 | new_G2872 | new_G2870 | new_G2871;
  assign G717 = ~new_G716;
  assign G820 = ~new_G819;
  assign new_G1046 = new_G2798 & G457;
  assign new_G1064 = new_G2794 & G468;
  assign new_G1071 = G422 & new_G2788;
  assign new_G1097 = new_G2784 & G435;
  assign new_G1111 = new_G2780 & G389;
  assign new_G1128 = new_G2776 & G400;
  assign new_G1145 = new_G2772 & G411;
  assign new_G1160 = new_G2767 & G374;
  assign new_G1301 = G457 & new_G2798;
  assign new_G1318 = G468 & new_G2794;
  assign new_G1324 = G422 & new_G2788;
  assign new_G1341 = G435 & new_G2784;
  assign new_G1359 = G389 & new_G2780;
  assign new_G1382 = G400 & new_G2776;
  assign new_G1404 = G411 & new_G2772;
  assign new_G1412 = G374 & new_G2767;
  assign new_G1704 = ~new_G3167;
  assign new_G1712 = ~new_G3165;
  assign new_G1724 = new_G3165;
  assign new_G1742 = new_G3161 & G479;
  assign new_G1749 = G490 & new_G3155;
  assign new_G1775 = new_G3151 & G503;
  assign new_G1806 = new_G3143 & G523;
  assign new_G1823 = new_G3139 & G534;
  assign new_G1829 = ~new_G3137;
  assign new_G1837 = new_G3137;
  assign new_G1958 = ~new_G3167;
  assign new_G1966 = ~new_G3165;
  assign new_G1978 = new_G3165;
  assign new_G1995 = G479 & new_G3161;
  assign new_G2001 = G490 & new_G3155;
  assign new_G2018 = G503 & new_G3151;
  assign new_G2059 = G523 & new_G3143;
  assign new_G2081 = G534 & new_G3139;
  assign new_G2089 = new_G3137;
  assign new_G2106 = ~new_G3137;
  assign new_G3170 = new_G3167;
  assign new_G3332 = ~new_G3331;
  assign new_G3339 = ~new_G3338;
  assign new_G5132 = ~new_G5126;
  assign new_G5184 = ~new_G5178;
  assign new_G3853 = ~new_G3852;
  assign new_G3874 = ~new_G3348;
  assign new_G4076 = new_G4056 & new_G2936 & new_G4037;
  assign new_G4116 = new_G2802;
  assign new_G4124 = new_G2798;
  assign new_G4132 = new_G2794;
  assign new_G4140 = new_G2788;
  assign new_G4148 = new_G2784;
  assign new_G4156 = new_G2780;
  assign new_G4164 = new_G2776;
  assign new_G4172 = new_G2772;
  assign new_G4180 = new_G2767;
  assign new_G4228 = ~G422 & ~new_G2788;
  assign new_G4279 = new_G2802;
  assign new_G4287 = new_G2798;
  assign new_G4295 = new_G2794;
  assign new_G4303 = new_G2784;
  assign new_G4311 = new_G2780;
  assign new_G4319 = new_G2776;
  assign new_G4327 = new_G2772;
  assign new_G4335 = new_G2788;
  assign new_G4343 = new_G2767;
  assign new_G4348 = ~G422 & ~new_G2788;
  assign new_G4464 = ~G374 & ~new_G2767;
  assign new_G4628 = new_G3161;
  assign new_G4636 = new_G3155;
  assign new_G4644 = new_G3151;
  assign new_G4660 = new_G3143;
  assign new_G4668 = new_G3139;
  assign new_G4716 = ~G490 & ~new_G3155;
  assign new_G4767 = new_G3161;
  assign new_G4775 = new_G3151;
  assign new_G4791 = new_G3143;
  assign new_G4799 = new_G3139;
  assign new_G4807 = new_G3155;
  assign new_G4812 = ~G490 & ~new_G3155;
  assign new_G5118 = new_G3139;
  assign new_G5121 = new_G3143;
  assign new_G5129 = new_G3137;
  assign new_G5134 = new_G3151;
  assign new_G5142 = new_G3161;
  assign new_G5145 = new_G3155;
  assign new_G5152 = new_G3167;
  assign new_G5155 = new_G3165;
  assign new_G5162 = new_G2788;
  assign new_G5165 = new_G2784;
  assign new_G5170 = new_G2798;
  assign new_G5173 = new_G2794;
  assign new_G5181 = new_G2802;
  assign new_G5186 = new_G2772;
  assign new_G5189 = new_G2767;
  assign new_G5196 = new_G2780;
  assign new_G5199 = new_G2776;
  assign new_G5214 = ~new_G5209 | ~new_G5212;
  assign new_G5215 = ~new_G5206 | ~new_G5213;
  assign new_G5329 = ~new_G5325;
  assign new_G5330 = ~new_G5325 | ~new_G5328;
  assign new_G2807 = ~new_G2942;
  assign new_G2808 = ~new_G2939;
  assign new_G2811 = ~new_G3021;
  assign new_G2812 = ~new_G3018;
  assign new_G2814 = ~new_G3012;
  assign new_G2626 = ~new_G2623;
  assign new_G2622 = ~new_G2619;
  assign new_G2618 = ~new_G2615;
  assign new_G2614 = ~new_G2611;
  assign new_G2720 = ~new_G2717;
  assign new_G2716 = ~new_G2713;
  assign new_G2712 = ~new_G2709;
  assign new_G2708 = ~new_G2705;
  assign G639 = new_G637 & new_G2827;
  assign G673 = new_G671 & new_G2827;
  assign G707 = new_G705 & new_G2827;
  assign G715 = new_G713 & new_G2827;
  assign new_G3731 = new_G3721 & new_G2945 & new_G3728;
  assign new_G4658 = ~new_G4652;
  assign new_G1777 = ~new_G4652 | ~new_G4659;
  assign new_G2019 = ~new_G4783 | ~new_G4786;
  assign new_G4787 = ~new_G4783;
  assign new_G3350 = new_G3332 & new_G3343;
  assign new_G3353 = new_G3339 & new_G3347;
  assign new_G5141 = ~new_G5137;
  assign new_G3513 = new_G3492 & new_G3428 & new_G3433;
  assign new_G3516 = new_G3496 & new_G3424 & new_G3437;
  assign new_G3517 = new_G3493 & new_G3437 & new_G3428;
  assign new_G3778 = new_G3765 & new_G2717 & new_G3745;
  assign new_G3781 = new_G3765 & new_G2713 & new_G3745;
  assign new_G3784 = new_G3765 & new_G2709 & new_G3745;
  assign new_G3787 = new_G3765 & new_G2705 & new_G3745;
  assign new_G3839 = new_G3823 & new_G3021 & new_G3803;
  assign new_G3842 = new_G3823 & new_G3018 & new_G3803;
  assign new_G5266 = ~new_G5260;
  assign new_G5267 = ~new_G5263;
  assign new_G5274 = ~new_G5268;
  assign new_G5275 = ~new_G5271;
  assign new_G5302 = ~new_G5296;
  assign new_G5303 = ~new_G5299;
  assign new_G5310 = ~new_G5304;
  assign new_G3891 = ~new_G5304 | ~new_G5311;
  assign new_G3937 = ~new_G3934;
  assign new_G3941 = ~new_G3938;
  assign new_G3955 = new_G3934 & new_G3906 & new_G3897;
  assign new_G3958 = new_G3938 & new_G3910 & new_G3901;
  assign new_G4009 = new_G3998 & new_G2623 & new_G3979;
  assign new_G4012 = new_G3998 & new_G2619 & new_G3979;
  assign new_G4015 = new_G3998 & new_G2615 & new_G3979;
  assign new_G4018 = new_G3998 & new_G2611 & new_G3979;
  assign new_G4067 = new_G4056 & new_G3012 & new_G4037;
  assign new_G4070 = new_G4056 & new_G2942 & new_G4037;
  assign new_G4073 = new_G4056 & new_G2939 & new_G4037;
  assign new_G4079 = new_G4056 & new_G2945 & new_G4037;
  assign new_G5239 = ~new_G5214 | ~new_G5215;
  assign new_G5282 = ~new_G5276;
  assign new_G5283 = ~new_G5279;
  assign new_G5293 = ~new_G5289;
  assign new_G5318 = ~new_G5312;
  assign new_G5319 = ~new_G5315;
  assign new_G5331 = ~new_G5322 | ~new_G5329;
  assign new_G5402 = ~new_G5396;
  assign new_G5405 = ~new_G5396 | ~new_G5403;
  assign new_G595 = new_G2810 & new_G2809 & new_G2807 & new_G2808;
  assign new_G596 = new_G2814 & new_G2813 & new_G2811 & new_G2812;
  assign new_G607 = new_G2614 & new_G2618 & new_G2626 & new_G2622;
  assign new_G608 = new_G2708 & new_G2712 & new_G2720 & new_G2716;
  assign new_G1845 = new_G1704 & new_G1724;
  assign new_G1846 = new_G1742 & new_G1712 & new_G1704;
  assign new_G2115 = new_G1958 & new_G1978;
  assign new_G2116 = new_G1995 & new_G1966 & new_G1958;
  assign new_G4122 = ~new_G4116;
  assign new_G1022 = ~new_G4116 | ~new_G4123;
  assign new_G4130 = ~new_G4124;
  assign new_G1033 = ~new_G4124 | ~new_G4131;
  assign new_G4138 = ~new_G4132;
  assign new_G1051 = ~new_G4132 | ~new_G4139;
  assign new_G4146 = ~new_G4140;
  assign new_G1079 = ~new_G4140 | ~new_G4147;
  assign new_G4154 = ~new_G4148;
  assign new_G1088 = ~new_G4148 | ~new_G4155;
  assign new_G4162 = ~new_G4156;
  assign new_G1099 = ~new_G4156 | ~new_G4163;
  assign new_G4170 = ~new_G4164;
  assign new_G1115 = ~new_G4164 | ~new_G4171;
  assign new_G4178 = ~new_G4172;
  assign new_G1133 = ~new_G4172 | ~new_G4179;
  assign new_G4186 = ~new_G4180;
  assign new_G1151 = ~new_G4180 | ~new_G4187;
  assign new_G4234 = ~new_G4228;
  assign new_G1276 = ~new_G4279 | ~new_G4282;
  assign new_G4283 = ~new_G4279;
  assign new_G1287 = ~new_G4287 | ~new_G4290;
  assign new_G4291 = ~new_G4287;
  assign new_G1305 = ~new_G4295 | ~new_G4298;
  assign new_G4299 = ~new_G4295;
  assign new_G1330 = ~new_G4303 | ~new_G4306;
  assign new_G4307 = ~new_G4303;
  assign new_G1342 = ~new_G4311 | ~new_G4314;
  assign new_G4315 = ~new_G4311;
  assign new_G1363 = ~new_G4319 | ~new_G4322;
  assign new_G4323 = ~new_G4319;
  assign new_G1388 = ~new_G4327 | ~new_G4330;
  assign new_G4331 = ~new_G4327;
  assign new_G1420 = ~new_G4335 | ~new_G4338;
  assign new_G4339 = ~new_G4335;
  assign new_G1428 = ~new_G4343 | ~new_G4346;
  assign new_G4347 = ~new_G4343;
  assign new_G4634 = ~new_G4628;
  assign new_G1729 = ~new_G4628 | ~new_G4635;
  assign new_G4642 = ~new_G4636;
  assign new_G1757 = ~new_G4636 | ~new_G4643;
  assign new_G4650 = ~new_G4644;
  assign new_G1766 = ~new_G4644 | ~new_G4651;
  assign new_G1776 = ~new_G4655 | ~new_G4658;
  assign new_G4666 = ~new_G4660;
  assign new_G1793 = ~new_G4660 | ~new_G4667;
  assign new_G4674 = ~new_G4668;
  assign new_G1811 = ~new_G4668 | ~new_G4675;
  assign new_G1849 = new_G1712 & new_G1742;
  assign new_G1852 = new_G1712 & new_G1742;
  assign new_G1875 = G54 & new_G1829;
  assign new_G4722 = ~new_G4716;
  assign new_G1982 = ~new_G4767 | ~new_G4770;
  assign new_G4771 = ~new_G4767;
  assign new_G2007 = ~new_G4775 | ~new_G4778;
  assign new_G4779 = ~new_G4775;
  assign new_G2020 = ~new_G4780 | ~new_G4787;
  assign new_G2040 = ~new_G4791 | ~new_G4794;
  assign new_G4795 = ~new_G4791;
  assign new_G2065 = ~new_G4799 | ~new_G4802;
  assign new_G4803 = ~new_G4799;
  assign new_G2097 = ~new_G4807 | ~new_G4810;
  assign new_G4811 = ~new_G4807;
  assign new_G2119 = new_G1966 & new_G1995;
  assign new_G2122 = new_G1966 & new_G1995;
  assign new_G5124 = ~new_G5118;
  assign new_G5125 = ~new_G5121;
  assign new_G3452 = ~new_G5129 | ~new_G5132;
  assign new_G5133 = ~new_G5129;
  assign new_G5140 = ~new_G5134;
  assign new_G3462 = ~new_G5134 | ~new_G5141;
  assign new_G5168 = ~new_G5162;
  assign new_G5169 = ~new_G5165;
  assign new_G5176 = ~new_G5170;
  assign new_G5177 = ~new_G5173;
  assign new_G3484 = ~new_G5181 | ~new_G5184;
  assign new_G5185 = ~new_G5181;
  assign new_G3515 = ~new_G3513 & ~new_G3514;
  assign new_G3518 = ~new_G3516 & ~new_G3517;
  assign new_G3857 = ~new_G3853;
  assign new_G3860 = ~new_G5263 | ~new_G5266;
  assign new_G3861 = ~new_G5260 | ~new_G5267;
  assign new_G3869 = ~new_G5271 | ~new_G5274;
  assign new_G3870 = ~new_G5268 | ~new_G5275;
  assign new_G3878 = ~new_G3874;
  assign new_G3881 = ~new_G5299 | ~new_G5302;
  assign new_G3882 = ~new_G5296 | ~new_G5303;
  assign new_G3890 = ~new_G5307 | ~new_G5310;
  assign new_G3954 = new_G3937 & new_G3901 & new_G3906;
  assign new_G3957 = new_G3941 & new_G3897 & new_G3910;
  assign new_G4021 = new_G3998 & new_G3353 & new_G3979;
  assign new_G4099 = ~new_G3170;
  assign new_G4236 = new_G1071;
  assign new_G4354 = ~new_G4348;
  assign new_G4406 = new_G1324;
  assign new_G4470 = ~new_G4464;
  assign new_G4552 = new_G1412;
  assign new_G4679 = new_G1829;
  assign new_G4687 = new_G1704;
  assign new_G4695 = new_G1704;
  assign new_G4703 = new_G1712;
  assign new_G4711 = new_G1712;
  assign new_G4724 = new_G1749;
  assign new_G4818 = ~new_G4812;
  assign new_G4855 = new_G1958;
  assign new_G4865 = new_G1966;
  assign new_G4870 = new_G2001;
  assign new_G4913 = new_G1958;
  assign new_G4923 = new_G1966;
  assign new_G4951 = new_G2106;
  assign new_G5006 = new_G2089;
  assign new_G5039 = new_G2106;
  assign new_G5148 = ~new_G5142;
  assign new_G5149 = ~new_G5145;
  assign new_G5158 = ~new_G5152;
  assign new_G5159 = ~new_G5155;
  assign new_G5192 = ~new_G5186;
  assign new_G5193 = ~new_G5189;
  assign new_G5202 = ~new_G5196;
  assign new_G5203 = ~new_G5199;
  assign new_G5284 = ~new_G5279 | ~new_G5282;
  assign new_G5285 = ~new_G5276 | ~new_G5283;
  assign new_G5320 = ~new_G5315 | ~new_G5318;
  assign new_G5321 = ~new_G5312 | ~new_G5319;
  assign new_G5386 = ~new_G5330 | ~new_G5331;
  assign new_G5404 = ~new_G5399 | ~new_G5402;
  assign G598 = new_G597 & new_G595 & new_G596;
  assign new_G609 = ~new_G3350;
  assign new_G1021 = ~new_G4119 | ~new_G4122;
  assign new_G1032 = ~new_G4127 | ~new_G4130;
  assign new_G1050 = ~new_G4135 | ~new_G4138;
  assign new_G1078 = ~new_G4143 | ~new_G4146;
  assign new_G1087 = ~new_G4151 | ~new_G4154;
  assign new_G1098 = ~new_G4159 | ~new_G4162;
  assign new_G1114 = ~new_G4167 | ~new_G4170;
  assign new_G1132 = ~new_G4175 | ~new_G4178;
  assign new_G1150 = ~new_G4183 | ~new_G4186;
  assign new_G1277 = ~new_G4276 | ~new_G4283;
  assign new_G1288 = ~new_G4284 | ~new_G4291;
  assign new_G1306 = ~new_G4292 | ~new_G4299;
  assign new_G1331 = ~new_G4300 | ~new_G4307;
  assign new_G1343 = ~new_G4308 | ~new_G4315;
  assign new_G1364 = ~new_G4316 | ~new_G4323;
  assign new_G1389 = ~new_G4324 | ~new_G4331;
  assign new_G1421 = ~new_G4332 | ~new_G4339;
  assign new_G1429 = ~new_G4340 | ~new_G4347;
  assign new_G1728 = ~new_G4631 | ~new_G4634;
  assign new_G1756 = ~new_G4639 | ~new_G4642;
  assign new_G1765 = ~new_G4647 | ~new_G4650;
  assign new_G1778 = ~new_G1776 | ~new_G1777;
  assign new_G1792 = ~new_G4663 | ~new_G4666;
  assign new_G1810 = ~new_G4671 | ~new_G4674;
  assign new_G1983 = ~new_G4764 | ~new_G4771;
  assign new_G2008 = ~new_G4772 | ~new_G4779;
  assign new_G2021 = ~new_G2019 | ~new_G2020;
  assign new_G2041 = ~new_G4788 | ~new_G4795;
  assign new_G2066 = ~new_G4796 | ~new_G4803;
  assign new_G2098 = ~new_G4804 | ~new_G4811;
  assign new_G3443 = ~new_G5121 | ~new_G5124;
  assign new_G3444 = ~new_G5118 | ~new_G5125;
  assign new_G3453 = ~new_G5126 | ~new_G5133;
  assign new_G3461 = ~new_G5137 | ~new_G5140;
  assign new_G3466 = ~new_G5165 | ~new_G5168;
  assign new_G3467 = ~new_G5162 | ~new_G5169;
  assign new_G3475 = ~new_G5173 | ~new_G5176;
  assign new_G3476 = ~new_G5170 | ~new_G5177;
  assign new_G3485 = ~new_G5178 | ~new_G5185;
  assign new_G5243 = ~new_G5239;
  assign new_G3862 = ~new_G3860 | ~new_G3861;
  assign new_G3871 = ~new_G3869 | ~new_G3870;
  assign new_G3883 = ~new_G3881 | ~new_G3882;
  assign new_G3892 = ~new_G3890 | ~new_G3891;
  assign new_G3956 = ~new_G3954 & ~new_G3955;
  assign new_G3959 = ~new_G3957 & ~new_G3958;
  assign new_G4756 = new_G1837 | new_G1875;
  assign new_G5150 = ~new_G5145 | ~new_G5148;
  assign new_G5151 = ~new_G5142 | ~new_G5149;
  assign new_G5160 = ~new_G5155 | ~new_G5158;
  assign new_G5161 = ~new_G5152 | ~new_G5159;
  assign new_G5194 = ~new_G5189 | ~new_G5192;
  assign new_G5195 = ~new_G5186 | ~new_G5193;
  assign new_G5204 = ~new_G5199 | ~new_G5202;
  assign new_G5205 = ~new_G5196 | ~new_G5203;
  assign new_G5236 = ~new_G3518 | ~new_G3515;
  assign new_G5286 = new_G3350;
  assign new_G5379 = ~new_G5284 | ~new_G5285;
  assign new_G5389 = ~new_G5320 | ~new_G5321;
  assign new_G5425 = ~new_G5404 | ~new_G5405;
  assign G610 = new_G609 & new_G607 & new_G608;
  assign new_G1023 = ~new_G1021 | ~new_G1022;
  assign new_G1034 = ~new_G1032 | ~new_G1033;
  assign new_G1052 = ~new_G1050 | ~new_G1051;
  assign new_G1080 = ~new_G1078 | ~new_G1079;
  assign new_G1089 = ~new_G1087 | ~new_G1088;
  assign new_G1100 = ~new_G1098 | ~new_G1099;
  assign new_G1116 = ~new_G1114 | ~new_G1115;
  assign new_G1134 = ~new_G1132 | ~new_G1133;
  assign new_G1152 = ~new_G1150 | ~new_G1151;
  assign new_G4242 = ~new_G4236;
  assign new_G1278 = ~new_G1276 | ~new_G1277;
  assign new_G1289 = ~new_G1287 | ~new_G1288;
  assign new_G1307 = ~new_G1305 | ~new_G1306;
  assign new_G1332 = ~new_G1330 | ~new_G1331;
  assign new_G1344 = ~new_G1342 | ~new_G1343;
  assign new_G1365 = ~new_G1363 | ~new_G1364;
  assign new_G1390 = ~new_G1388 | ~new_G1389;
  assign new_G1422 = ~new_G1420 | ~new_G1421;
  assign new_G1430 = ~new_G1428 | ~new_G1429;
  assign new_G1730 = ~new_G1728 | ~new_G1729;
  assign new_G1758 = ~new_G1756 | ~new_G1757;
  assign new_G1767 = ~new_G1765 | ~new_G1766;
  assign new_G1794 = ~new_G1792 | ~new_G1793;
  assign new_G1812 = ~new_G1810 | ~new_G1811;
  assign new_G1876 = ~new_G4679 | ~new_G4682;
  assign new_G4683 = ~new_G4679;
  assign new_G4691 = ~new_G4687;
  assign new_G4699 = ~new_G4695;
  assign new_G4707 = ~new_G4703;
  assign new_G4715 = ~new_G4711;
  assign new_G4730 = ~new_G4724;
  assign new_G1984 = ~new_G1982 | ~new_G1983;
  assign new_G2009 = ~new_G2007 | ~new_G2008;
  assign new_G2042 = ~new_G2040 | ~new_G2041;
  assign new_G2067 = ~new_G2065 | ~new_G2066;
  assign new_G2099 = ~new_G2097 | ~new_G2098;
  assign new_G4869 = ~new_G4865;
  assign new_G4927 = ~new_G4923;
  assign new_G3445 = ~new_G3443 | ~new_G3444;
  assign new_G3454 = ~new_G3452 | ~new_G3453;
  assign new_G3463 = ~new_G3461 | ~new_G3462;
  assign new_G3468 = ~new_G3466 | ~new_G3467;
  assign new_G3477 = ~new_G3475 | ~new_G3476;
  assign new_G3486 = ~new_G3484 | ~new_G3485;
  assign new_G4103 = new_G4099 & new_G3170;
  assign new_G4412 = ~new_G4406;
  assign new_G4558 = ~new_G4552;
  assign new_G4859 = ~new_G4855;
  assign new_G4876 = ~new_G4870;
  assign new_G4917 = ~new_G4913;
  assign new_G4955 = ~new_G4951;
  assign new_G5012 = ~new_G5006;
  assign new_G5043 = ~new_G5039;
  assign new_G5216 = ~new_G5160 | ~new_G5161;
  assign new_G5219 = ~new_G5150 | ~new_G5151;
  assign new_G5226 = ~new_G5204 | ~new_G5205;
  assign new_G5229 = ~new_G5194 | ~new_G5195;
  assign new_G5392 = ~new_G5386;
  assign new_G5422 = ~new_G3959 | ~new_G3956;
  assign new_G1866 = new_G1778 & new_G1806;
  assign new_G1877 = ~new_G4676 | ~new_G4683;
  assign new_G4762 = ~new_G4756;
  assign new_G2142 = new_G2021 & new_G2059;
  assign new_G2146 = new_G2021 & new_G2059;
  assign new_G5242 = ~new_G5236;
  assign new_G3532 = ~new_G5236 | ~new_G5243;
  assign new_G3866 = ~new_G3862;
  assign new_G3887 = ~new_G3883;
  assign new_G3918 = new_G3871;
  assign new_G3922 = new_G3871;
  assign new_G3926 = new_G3892;
  assign new_G3930 = new_G3892;
  assign new_G5429 = ~new_G5425;
  assign new_G4104 = new_G4099 | new_G4103;
  assign new_G4743 = new_G1778;
  assign new_G4991 = new_G2021;
  assign new_G5001 = new_G2021;
  assign new_G5292 = ~new_G5286;
  assign new_G5295 = ~new_G5286 | ~new_G5293;
  assign new_G5383 = ~new_G5379;
  assign new_G5393 = ~new_G5389;
  assign new_G5394 = ~new_G5389 | ~new_G5392;
  assign new_G1439 = new_G1278 & new_G1301;
  assign new_G1440 = new_G1318 & new_G1289 & new_G1278;
  assign new_G1441 = new_G1289 & new_G1324 & new_G1307 & new_G1278;
  assign new_G1847 = new_G1712 & new_G1749 & new_G1730 & new_G1704;
  assign new_G1168 = new_G1023 & new_G1046;
  assign new_G1169 = new_G1064 & new_G1034 & new_G1023;
  assign new_G1170 = new_G1034 & new_G1071 & new_G1052 & new_G1023;
  assign new_G2117 = new_G1966 & new_G2001 & new_G1984 & new_G1958;
  assign new_G1086 = ~new_G1080;
  assign new_G1166 = new_G1023 & new_G1052 & new_G1034 & new_G1080;
  assign new_G1171 = new_G1034 & new_G1064;
  assign new_G1172 = new_G1034 & new_G1052 & new_G1071;
  assign new_G1173 = new_G1034 & new_G1080 & new_G1052;
  assign new_G1174 = new_G1034 & new_G1064;
  assign new_G1175 = new_G1034 & new_G1071 & new_G1052;
  assign new_G1176 = new_G1052 & new_G1071;
  assign new_G1177 = new_G1080 & new_G1052;
  assign new_G1178 = new_G1052 & new_G1071;
  assign new_G1179 = new_G1134 & new_G1089 & new_G1116 & new_G1100 & new_G1152;
  assign new_G1181 = new_G1089 & new_G1111;
  assign new_G1182 = new_G1128 & new_G1100 & new_G1089;
  assign new_G1183 = new_G1100 & new_G1145 & new_G1116 & new_G1089;
  assign new_G1184 = new_G1100 & new_G1160 & new_G1089 & new_G1134 & new_G1116;
  assign new_G1188 = new_G1100 & new_G1128;
  assign new_G1189 = new_G1100 & new_G1116 & new_G1145;
  assign new_G1190 = new_G1100 & new_G1160 & new_G1134 & new_G1116;
  assign new_G1191 = new_G1100 & new_G1134 & new_G1116 & G4 & new_G1152;
  assign new_G1192 = new_G1145 & new_G1116;
  assign new_G1193 = new_G1160 & new_G1134 & new_G1116;
  assign new_G1194 = new_G1134 & new_G1116 & G4 & new_G1152;
  assign new_G1195 = new_G1134 & new_G1160;
  assign new_G1196 = new_G1134 & G4 & new_G1152;
  assign new_G1197 = G4 & new_G1152;
  assign new_G1437 = new_G1278 & new_G1289 & new_G1422 & new_G1307;
  assign new_G1442 = new_G1289 & new_G1318;
  assign new_G1443 = new_G1289 & new_G1307 & new_G1324;
  assign new_G1444 = new_G1289 & new_G1422 & new_G1307;
  assign new_G1445 = new_G1289 & new_G1318;
  assign new_G1446 = new_G1289 & new_G1307 & new_G1324;
  assign new_G1447 = new_G1307 & new_G1324;
  assign new_G1451 = new_G1332 & new_G1344 & new_G1365 & new_G1430 & new_G1390;
  assign new_G1454 = new_G1332 & new_G1359;
  assign new_G1455 = new_G1382 & new_G1344 & new_G1332;
  assign new_G1456 = new_G1344 & new_G1404 & new_G1365 & new_G1332;
  assign new_G1457 = new_G1344 & new_G1412 & new_G1332 & new_G1390 & new_G1365;
  assign new_G1465 = new_G1344 & new_G1382;
  assign new_G1466 = new_G1344 & new_G1365 & new_G1404;
  assign new_G1467 = new_G1344 & new_G1412 & new_G1390 & new_G1365;
  assign new_G1468 = new_G1390 & new_G1344 & new_G1430 & new_G1365;
  assign new_G1469 = new_G1344 & new_G1382;
  assign new_G1470 = new_G1344 & new_G1365 & new_G1404;
  assign new_G1471 = new_G1344 & new_G1412 & new_G1390 & new_G1365;
  assign new_G1472 = new_G1365 & new_G1404;
  assign new_G1473 = new_G1412 & new_G1390 & new_G1365;
  assign new_G1474 = new_G1390 & new_G1430 & new_G1365;
  assign new_G1475 = new_G1365 & new_G1404;
  assign new_G1476 = new_G1412 & new_G1390 & new_G1365;
  assign new_G1477 = new_G1390 & new_G1412;
  assign new_G1481 = new_G1422 & new_G1307;
  assign new_G1482 = new_G1430 & new_G1390;
  assign new_G1764 = ~new_G1758;
  assign new_G1843 = new_G1704 & new_G1730 & new_G1712 & new_G1758;
  assign new_G1850 = new_G1712 & new_G1730 & new_G1749;
  assign new_G1851 = new_G1712 & new_G1758 & new_G1730;
  assign new_G1853 = new_G1712 & new_G1749 & new_G1730;
  assign new_G1854 = new_G1730 & new_G1749;
  assign new_G1855 = new_G1758 & new_G1730;
  assign new_G1856 = new_G1730 & new_G1749;
  assign new_G1857 = new_G1812 & new_G1767 & new_G1794 & new_G1778 & new_G1829;
  assign new_G1859 = new_G1767 & new_G1789;
  assign new_G1860 = new_G1806 & new_G1778 & new_G1767;
  assign new_G1861 = new_G1778 & new_G1823 & new_G1794 & new_G1767;
  assign new_G1862 = new_G1778 & new_G1837 & new_G1767 & new_G1812 & new_G1794;
  assign new_G1867 = new_G1778 & new_G1794 & new_G1823;
  assign new_G1868 = new_G1778 & new_G1837 & new_G1812 & new_G1794;
  assign new_G1869 = new_G1778 & new_G1812 & new_G1794 & G54 & new_G1829;
  assign new_G1870 = new_G1823 & new_G1794;
  assign new_G1871 = new_G1837 & new_G1812 & new_G1794;
  assign new_G1872 = new_G1812 & new_G1794 & G54 & new_G1829;
  assign new_G1873 = new_G1812 & new_G1837;
  assign new_G1874 = new_G1812 & G54 & new_G1829;
  assign new_G1878 = ~new_G1876 | ~new_G1877;
  assign new_G2113 = new_G1958 & new_G1966 & new_G2099 & new_G1984;
  assign new_G2120 = new_G1966 & new_G1984 & new_G2001;
  assign new_G2121 = new_G1966 & new_G2099 & new_G1984;
  assign new_G2123 = new_G1966 & new_G1984 & new_G2001;
  assign new_G2124 = new_G1984 & new_G2001;
  assign new_G2128 = new_G2009 & new_G2021 & new_G2042 & new_G2106 & new_G2067;
  assign new_G2131 = new_G2009 & new_G2036;
  assign new_G2132 = new_G2059 & new_G2021 & new_G2009;
  assign new_G2133 = new_G2021 & new_G2081 & new_G2042 & new_G2009;
  assign new_G2134 = new_G2021 & new_G2089 & new_G2009 & new_G2067 & new_G2042;
  assign new_G2143 = new_G2021 & new_G2042 & new_G2081;
  assign new_G2144 = new_G2021 & new_G2089 & new_G2067 & new_G2042;
  assign new_G2145 = new_G2067 & new_G2021 & new_G2106 & new_G2042;
  assign new_G2147 = new_G2021 & new_G2042 & new_G2081;
  assign new_G2148 = new_G2021 & new_G2089 & new_G2067 & new_G2042;
  assign new_G2149 = new_G2042 & new_G2081;
  assign new_G2150 = new_G2089 & new_G2067 & new_G2042;
  assign new_G2151 = new_G2067 & new_G2106 & new_G2042;
  assign new_G2152 = new_G2042 & new_G2081;
  assign new_G2153 = new_G2089 & new_G2067 & new_G2042;
  assign new_G2154 = new_G2067 & new_G2089;
  assign new_G2158 = new_G2099 & new_G1984;
  assign new_G2159 = new_G2106 & new_G2067;
  assign new_G3449 = ~new_G3445;
  assign new_G3458 = ~new_G3454;
  assign new_G3472 = ~new_G3468;
  assign new_G3481 = ~new_G3477;
  assign new_G3497 = new_G3463;
  assign new_G3501 = new_G3463;
  assign new_G3505 = new_G3486;
  assign new_G3509 = new_G3486;
  assign new_G3531 = ~new_G5239 | ~new_G5242;
  assign new_G5428 = ~new_G5422;
  assign new_G3967 = ~new_G5422 | ~new_G5429;
  assign new_G4191 = new_G1152;
  assign new_G4199 = new_G1023;
  assign new_G4207 = new_G1023;
  assign new_G4215 = new_G1034;
  assign new_G4223 = new_G1034;
  assign new_G4231 = new_G1052;
  assign new_G4239 = new_G1052;
  assign new_G4247 = new_G1089;
  assign new_G4255 = new_G1100;
  assign new_G4263 = new_G1116;
  assign new_G4271 = new_G1134;
  assign new_G4371 = new_G1422;
  assign new_G4381 = new_G1307;
  assign new_G4391 = new_G1278;
  assign new_G4401 = new_G1289;
  assign new_G4429 = new_G1422;
  assign new_G4439 = new_G1307;
  assign new_G4449 = new_G1278;
  assign new_G4459 = new_G1289;
  assign new_G4497 = new_G1430;
  assign new_G4507 = new_G1390;
  assign new_G4517 = new_G1332;
  assign new_G4527 = new_G1365;
  assign new_G4537 = new_G1344;
  assign new_G4547 = new_G1344;
  assign new_G4585 = new_G1430;
  assign new_G4595 = new_G1390;
  assign new_G4605 = new_G1332;
  assign new_G4615 = new_G1365;
  assign new_G4719 = new_G1730;
  assign new_G4727 = new_G1730;
  assign new_G4735 = new_G1767;
  assign new_G4751 = new_G1794;
  assign new_G4759 = new_G1812;
  assign new_G4835 = new_G2099;
  assign new_G4845 = new_G1984;
  assign new_G4893 = new_G2099;
  assign new_G4903 = new_G1984;
  assign new_G4961 = new_G2067;
  assign new_G4971 = new_G2009;
  assign new_G4981 = new_G2042;
  assign new_G5049 = new_G2067;
  assign new_G5059 = new_G2009;
  assign new_G5069 = new_G2042;
  assign new_G5222 = ~new_G5216;
  assign new_G5223 = ~new_G5219;
  assign new_G5232 = ~new_G5226;
  assign new_G5233 = ~new_G5229;
  assign new_G5294 = ~new_G5289 | ~new_G5292;
  assign new_G5395 = ~new_G5386 | ~new_G5393;
  assign new_G589 = new_G1441 | new_G1440 | new_G1286 | new_G1439;
  assign new_G616 = new_G1847 | new_G1846 | new_G3167 | new_G1845;
  assign new_G619 = new_G1170 | new_G1169 | new_G1031 | new_G1168;
  assign new_G627 = new_G2117 | new_G2116 | new_G3167 | new_G2115;
  assign new_G1185 = new_G1184 | new_G1183 | new_G1182 | new_G1097 | new_G1181;
  assign new_G1448 = new_G1318 | new_G1447;
  assign new_G1458 = new_G1457 | new_G1456 | new_G1455 | new_G1341 | new_G1454;
  assign new_G1478 = new_G1404 | new_G1477;
  assign new_G1863 = new_G1862 | new_G1861 | new_G1860 | new_G1775 | new_G1859;
  assign new_G4747 = ~new_G4743;
  assign new_G2125 = new_G1995 | new_G2124;
  assign new_G2135 = new_G2134 | new_G2133 | new_G2132 | new_G2018 | new_G2131;
  assign new_G2155 = new_G2081 | new_G2154;
  assign new_G4995 = ~new_G4991;
  assign new_G5005 = ~new_G5001;
  assign new_G3533 = ~new_G3531 | ~new_G3532;
  assign new_G3921 = ~new_G3918;
  assign new_G3925 = ~new_G3922;
  assign new_G3929 = ~new_G3926;
  assign new_G3933 = ~new_G3930;
  assign new_G3943 = new_G3918 & new_G3862 & new_G3853;
  assign new_G3946 = new_G3922 & new_G3866 & new_G3857;
  assign new_G3949 = new_G3926 & new_G3883 & new_G3874;
  assign new_G3952 = new_G3930 & new_G3887 & new_G3878;
  assign new_G3966 = ~new_G5425 | ~new_G5428;
  assign new_G4107 = ~new_G4104 | ~G132;
  assign new_G4196 = new_G1173 | new_G1172 | new_G1046 | new_G1171;
  assign new_G4204 = ~new_G1175 & ~new_G1046 & ~new_G1174;
  assign new_G4212 = new_G1177 | new_G1064 | new_G1176;
  assign new_G4220 = ~new_G1064 & ~new_G1178;
  assign new_G4244 = new_G1191 | new_G1190 | new_G1189 | new_G1111 | new_G1188;
  assign new_G4252 = new_G1194 | new_G1193 | new_G1128 | new_G1192;
  assign new_G4260 = new_G1196 | new_G1145 | new_G1195;
  assign new_G4268 = new_G1160 | new_G1197;
  assign new_G4361 = new_G1444 | new_G1443 | new_G1301 | new_G1442;
  assign new_G4419 = ~new_G1446 & ~new_G1301 & ~new_G1445;
  assign new_G4467 = new_G1474 | new_G1473 | new_G1382 | new_G1472;
  assign new_G4487 = new_G1468 | new_G1467 | new_G1466 | new_G1359 | new_G1465;
  assign new_G4555 = ~new_G1476 & ~new_G1382 & ~new_G1475;
  assign new_G4575 = ~new_G1471 & ~new_G1470 & ~new_G1359 & ~new_G1469;
  assign new_G4684 = new_G1851 | new_G1850 | new_G1724 | new_G1849;
  assign new_G4692 = ~new_G1853 & ~new_G1724 & ~new_G1852;
  assign new_G4700 = new_G1855 | new_G1742 | new_G1854;
  assign new_G4708 = ~new_G1742 & ~new_G1856;
  assign new_G4732 = new_G1869 | new_G1868 | new_G1867 | new_G1789 | new_G1866;
  assign new_G4740 = new_G1872 | new_G1871 | new_G1806 | new_G1870;
  assign new_G4748 = new_G1874 | new_G1823 | new_G1873;
  assign new_G4825 = new_G2121 | new_G2120 | new_G1978 | new_G2119;
  assign new_G4883 = ~new_G2123 & ~new_G1978 & ~new_G2122;
  assign new_G4928 = new_G2151 | new_G2150 | new_G2059 | new_G2149;
  assign new_G4941 = new_G2145 | new_G2144 | new_G2143 | new_G2036 | new_G2142;
  assign new_G5009 = ~new_G2153 & ~new_G2059 & ~new_G2152;
  assign new_G5029 = ~new_G2148 & ~new_G2147 & ~new_G2036 & ~new_G2146;
  assign new_G5224 = ~new_G5219 | ~new_G5222;
  assign new_G5225 = ~new_G5216 | ~new_G5223;
  assign new_G5234 = ~new_G5229 | ~new_G5232;
  assign new_G5235 = ~new_G5226 | ~new_G5233;
  assign new_G5376 = ~new_G5294 | ~new_G5295;
  assign new_G5417 = ~new_G5394 | ~new_G5395;
  assign new_G576 = ~new_G1878;
  assign G588 = new_G1437 & new_G1451;
  assign G615 = new_G1843 & new_G1857;
  assign G626 = new_G2113 & new_G2128;
  assign G632 = new_G1166 & new_G1179;
  assign new_G1198 = ~new_G4191 | ~new_G4194;
  assign new_G4195 = ~new_G4191;
  assign new_G4203 = ~new_G4199;
  assign new_G4211 = ~new_G4207;
  assign new_G4219 = ~new_G4215;
  assign new_G4227 = ~new_G4223;
  assign new_G1217 = ~new_G4231 | ~new_G4234;
  assign new_G4235 = ~new_G4231;
  assign new_G1221 = ~new_G4239 | ~new_G4242;
  assign new_G4243 = ~new_G4239;
  assign new_G1224 = new_G1179 & G4;
  assign new_G4251 = ~new_G4247;
  assign new_G4259 = ~new_G4255;
  assign new_G4267 = ~new_G4263;
  assign new_G4275 = ~new_G4271;
  assign new_G1453 = ~new_G1451;
  assign new_G4405 = ~new_G4401;
  assign new_G4463 = ~new_G4459;
  assign new_G4541 = ~new_G4537;
  assign new_G4551 = ~new_G4547;
  assign new_G1895 = ~new_G4719 | ~new_G4722;
  assign new_G4723 = ~new_G4719;
  assign new_G1899 = ~new_G4727 | ~new_G4730;
  assign new_G4731 = ~new_G4727;
  assign new_G1902 = new_G1857 & G54;
  assign new_G4739 = ~new_G4735;
  assign new_G4755 = ~new_G4751;
  assign new_G1929 = ~new_G4759 | ~new_G4762;
  assign new_G4763 = ~new_G4759;
  assign new_G2130 = ~new_G2128;
  assign new_G3500 = ~new_G3497;
  assign new_G3504 = ~new_G3501;
  assign new_G3508 = ~new_G3505;
  assign new_G3512 = ~new_G3509;
  assign new_G3520 = new_G3497 & new_G3454 & new_G3445;
  assign new_G3523 = new_G3501 & new_G3458 & new_G3449;
  assign new_G3526 = new_G3505 & new_G3477 & new_G3468;
  assign new_G3529 = new_G3509 & new_G3481 & new_G3472;
  assign G1002 = new_G3533;
  assign new_G3837 = new_G3823 & new_G1878 & new_G3795;
  assign new_G3942 = new_G3921 & new_G3857 & new_G3862;
  assign new_G3945 = new_G3925 & new_G3853 & new_G3866;
  assign new_G3948 = new_G3929 & new_G3878 & new_G3883;
  assign new_G3951 = new_G3933 & new_G3874 & new_G3887;
  assign new_G3968 = ~new_G3966 | ~new_G3967;
  assign new_G4375 = ~new_G4371;
  assign new_G4385 = ~new_G4381;
  assign new_G4395 = ~new_G4391;
  assign new_G4433 = ~new_G4429;
  assign new_G4443 = ~new_G4439;
  assign new_G4453 = ~new_G4449;
  assign new_G4501 = ~new_G4497;
  assign new_G4511 = ~new_G4507;
  assign new_G4521 = ~new_G4517;
  assign new_G4531 = ~new_G4527;
  assign new_G4619 = ~new_G4615;
  assign new_G4589 = ~new_G4585;
  assign new_G4599 = ~new_G4595;
  assign new_G4609 = ~new_G4605;
  assign new_G4839 = ~new_G4835;
  assign new_G4849 = ~new_G4845;
  assign new_G4897 = ~new_G4893;
  assign new_G4907 = ~new_G4903;
  assign new_G4965 = ~new_G4961;
  assign new_G4975 = ~new_G4971;
  assign new_G4985 = ~new_G4981;
  assign new_G5073 = ~new_G5069;
  assign new_G5053 = ~new_G5049;
  assign new_G5063 = ~new_G5059;
  assign new_G5247 = ~new_G5224 | ~new_G5225;
  assign new_G5255 = ~new_G5234 | ~new_G5235;
  assign new_G590 = new_G1437 & new_G1458;
  assign new_G617 = new_G1863 & new_G1843;
  assign new_G620 = new_G1185 & new_G1166;
  assign new_G628 = new_G2113 & new_G2135;
  assign new_G3535 = ~new_G3533;
  assign new_G1199 = ~new_G4188 | ~new_G4195;
  assign new_G4202 = ~new_G4196;
  assign new_G1204 = ~new_G4196 | ~new_G4203;
  assign new_G4210 = ~new_G4204;
  assign new_G1207 = ~new_G4204 | ~new_G4211;
  assign new_G4218 = ~new_G4212;
  assign new_G1211 = ~new_G4212 | ~new_G4219;
  assign new_G4226 = ~new_G4220;
  assign new_G1214 = ~new_G4220 | ~new_G4227;
  assign new_G1218 = ~new_G4228 | ~new_G4235;
  assign new_G1222 = ~new_G4236 | ~new_G4243;
  assign new_G1225 = new_G1185 | new_G1224;
  assign new_G4250 = ~new_G4244;
  assign new_G1237 = ~new_G4244 | ~new_G4251;
  assign new_G4258 = ~new_G4252;
  assign new_G1242 = ~new_G4252 | ~new_G4259;
  assign new_G4266 = ~new_G4260;
  assign new_G1247 = ~new_G4260 | ~new_G4267;
  assign new_G4274 = ~new_G4268;
  assign new_G1252 = ~new_G4268 | ~new_G4275;
  assign new_G1462 = ~new_G1458;
  assign new_G4690 = ~new_G4684;
  assign new_G1882 = ~new_G4684 | ~new_G4691;
  assign new_G4698 = ~new_G4692;
  assign new_G1885 = ~new_G4692 | ~new_G4699;
  assign new_G4706 = ~new_G4700;
  assign new_G1889 = ~new_G4700 | ~new_G4707;
  assign new_G4714 = ~new_G4708;
  assign new_G1892 = ~new_G4708 | ~new_G4715;
  assign new_G1896 = ~new_G4716 | ~new_G4723;
  assign new_G1900 = ~new_G4724 | ~new_G4731;
  assign new_G1903 = new_G1863 | new_G1902;
  assign new_G4738 = ~new_G4732;
  assign new_G1915 = ~new_G4732 | ~new_G4739;
  assign new_G4746 = ~new_G4740;
  assign new_G1920 = ~new_G4740 | ~new_G4747;
  assign new_G4754 = ~new_G4748;
  assign new_G1925 = ~new_G4748 | ~new_G4755;
  assign new_G1930 = ~new_G4756 | ~new_G4763;
  assign new_G2139 = ~new_G2135;
  assign new_G3519 = new_G3500 & new_G3449 & new_G3454;
  assign new_G3522 = new_G3504 & new_G3445 & new_G3458;
  assign new_G3525 = new_G3508 & new_G3472 & new_G3477;
  assign new_G3528 = new_G3512 & new_G3468 & new_G3481;
  assign new_G3848 = new_G3838 | new_G3836 | new_G3837;
  assign new_G3944 = ~new_G3942 & ~new_G3943;
  assign new_G3947 = ~new_G3945 & ~new_G3946;
  assign new_G3950 = ~new_G3948 & ~new_G3949;
  assign new_G3953 = ~new_G3951 & ~new_G3952;
  assign new_G5421 = ~new_G5417;
  assign G1004 = new_G3968;
  assign new_G4111 = new_G4104 & new_G4107;
  assign new_G4112 = new_G4107 & G132;
  assign new_G4351 = new_G1448 | new_G1481;
  assign new_G4365 = ~new_G4361;
  assign new_G4409 = ~new_G1448;
  assign new_G4423 = ~new_G4419;
  assign new_G4471 = ~new_G4467;
  assign new_G4472 = ~new_G4467 | ~new_G4470;
  assign new_G4477 = new_G1478 | new_G1482;
  assign new_G4491 = ~new_G4487;
  assign new_G4559 = ~new_G4555;
  assign new_G4560 = ~new_G4555 | ~new_G4558;
  assign new_G4565 = ~new_G1478;
  assign new_G4579 = ~new_G4575;
  assign new_G4815 = new_G2125 | new_G2158;
  assign new_G4829 = ~new_G4825;
  assign new_G4873 = ~new_G2125;
  assign new_G4887 = ~new_G4883;
  assign new_G4931 = new_G2155 | new_G2159;
  assign new_G4934 = ~new_G4928;
  assign new_G4945 = ~new_G4941;
  assign new_G5013 = ~new_G5009;
  assign new_G5014 = ~new_G5009 | ~new_G5012;
  assign new_G5019 = ~new_G2155;
  assign new_G5033 = ~new_G5029;
  assign new_G5382 = ~new_G5376;
  assign new_G5385 = ~new_G5376 | ~new_G5383;
  assign G591 = new_G589 | new_G590;
  assign G618 = new_G616 | new_G617;
  assign G621 = new_G619 | new_G620;
  assign G629 = new_G627 | new_G628;
  assign new_G3970 = ~new_G3968;
  assign new_G1200 = ~new_G1198 | ~new_G1199;
  assign new_G1203 = ~new_G4199 | ~new_G4202;
  assign new_G1206 = ~new_G4207 | ~new_G4210;
  assign new_G1210 = ~new_G4215 | ~new_G4218;
  assign new_G1213 = ~new_G4223 | ~new_G4226;
  assign new_G1219 = ~new_G1217 | ~new_G1218;
  assign new_G1223 = ~new_G1221 | ~new_G1222;
  assign new_G1236 = ~new_G4247 | ~new_G4250;
  assign new_G1241 = ~new_G4255 | ~new_G4258;
  assign new_G1246 = ~new_G4263 | ~new_G4266;
  assign new_G1251 = ~new_G4271 | ~new_G4274;
  assign new_G1881 = ~new_G4687 | ~new_G4690;
  assign new_G1884 = ~new_G4695 | ~new_G4698;
  assign new_G1888 = ~new_G4703 | ~new_G4706;
  assign new_G1891 = ~new_G4711 | ~new_G4714;
  assign new_G1897 = ~new_G1895 | ~new_G1896;
  assign new_G1901 = ~new_G1899 | ~new_G1900;
  assign new_G1914 = ~new_G4735 | ~new_G4738;
  assign new_G1919 = ~new_G4743 | ~new_G4746;
  assign new_G1924 = ~new_G4751 | ~new_G4754;
  assign new_G1931 = ~new_G1929 | ~new_G1930;
  assign new_G3521 = ~new_G3519 & ~new_G3520;
  assign new_G3524 = ~new_G3522 & ~new_G3523;
  assign new_G3527 = ~new_G3525 & ~new_G3526;
  assign new_G3530 = ~new_G3528 & ~new_G3529;
  assign new_G5251 = ~new_G5247;
  assign new_G5259 = ~new_G5255;
  assign new_G4113 = new_G4111 | new_G4112;
  assign new_G4473 = ~new_G4464 | ~new_G4471;
  assign new_G4561 = ~new_G4552 | ~new_G4559;
  assign new_G5015 = ~new_G5006 | ~new_G5013;
  assign new_G5384 = ~new_G5379 | ~new_G5382;
  assign new_G5406 = ~new_G3947 | ~new_G3944;
  assign new_G5414 = ~new_G3953 | ~new_G3950;
  assign new_G1664 = new_G1645 & new_G3848 & new_G1621;
  assign new_G2335 = new_G2316 & new_G3848 & new_G2293;
  assign new_G718 = new_G2454 & new_G3848 & new_G2430;
  assign G822 = ~new_G3848;
  assign new_G855 = new_G2512 & new_G3848 & new_G2488;
  assign new_G1205 = ~new_G1203 | ~new_G1204;
  assign new_G1208 = ~new_G1206 | ~new_G1207;
  assign new_G1212 = ~new_G1210 | ~new_G1211;
  assign new_G1215 = ~new_G1213 | ~new_G1214;
  assign new_G1220 = ~new_G1219;
  assign new_G1231 = ~new_G1225;
  assign new_G1238 = ~new_G1236 | ~new_G1237;
  assign new_G1243 = ~new_G1241 | ~new_G1242;
  assign new_G1248 = ~new_G1246 | ~new_G1247;
  assign new_G1253 = ~new_G1251 | ~new_G1252;
  assign new_G1272 = new_G1225 & new_G1086;
  assign new_G1483 = new_G1462 & new_G1453;
  assign new_G1883 = ~new_G1881 | ~new_G1882;
  assign new_G1886 = ~new_G1884 | ~new_G1885;
  assign new_G1890 = ~new_G1888 | ~new_G1889;
  assign new_G1893 = ~new_G1891 | ~new_G1892;
  assign new_G1898 = ~new_G1897;
  assign new_G1909 = ~new_G1903;
  assign new_G1916 = ~new_G1914 | ~new_G1915;
  assign new_G1921 = ~new_G1919 | ~new_G1920;
  assign new_G1926 = ~new_G1924 | ~new_G1925;
  assign new_G1953 = new_G1903 & new_G1764;
  assign new_G2160 = new_G2139 & new_G2130;
  assign new_G4355 = ~new_G4351;
  assign new_G4356 = ~new_G4351 | ~new_G4354;
  assign new_G4413 = ~new_G4409;
  assign new_G4414 = ~new_G4409 | ~new_G4412;
  assign new_G4474 = ~new_G4472 | ~new_G4473;
  assign new_G4481 = ~new_G4477;
  assign new_G4562 = ~new_G4560 | ~new_G4561;
  assign new_G4569 = ~new_G4565;
  assign new_G4819 = ~new_G4815;
  assign new_G4820 = ~new_G4815 | ~new_G4818;
  assign new_G4877 = ~new_G4873;
  assign new_G4878 = ~new_G4873 | ~new_G4876;
  assign new_G4935 = ~new_G4931;
  assign new_G4936 = ~new_G4931 | ~new_G4934;
  assign new_G5016 = ~new_G5014 | ~new_G5015;
  assign new_G5023 = ~new_G5019;
  assign new_G5244 = ~new_G3524 | ~new_G3521;
  assign new_G5252 = ~new_G3530 | ~new_G3527;
  assign new_G5409 = ~new_G5384 | ~new_G5385;
  assign new_G566 = ~new_G1200;
  assign new_G577 = ~new_G1931;
  assign new_G3733 = new_G3721 & new_G4113 & G3724;
  assign new_G1209 = ~new_G1208;
  assign new_G1216 = ~new_G1215;
  assign new_G1257 = new_G1225 & new_G1205;
  assign new_G1262 = new_G1225 & new_G1212;
  assign new_G1267 = new_G1225 & new_G1220;
  assign new_G1887 = ~new_G1886;
  assign new_G1894 = ~new_G1893;
  assign new_G1935 = new_G1903 & new_G1883;
  assign new_G1943 = new_G1903 & new_G1890;
  assign new_G1948 = new_G1903 & new_G1898;
  assign new_G3779 = new_G3765 & new_G1200 & new_G3737;
  assign new_G3840 = new_G3823 & new_G1931 & new_G3795;
  assign new_G5412 = ~new_G5406;
  assign new_G5420 = ~new_G5414;
  assign new_G3964 = ~new_G5414 | ~new_G5421;
  assign new_G4357 = ~new_G4348 | ~new_G4355;
  assign new_G4415 = ~new_G4406 | ~new_G4413;
  assign new_G4821 = ~new_G4812 | ~new_G4819;
  assign new_G4879 = ~new_G4870 | ~new_G4877;
  assign new_G4937 = ~new_G4928 | ~new_G4935;
  assign new_G567 = ~new_G1253;
  assign new_G568 = ~new_G1248;
  assign new_G569 = ~new_G1243;
  assign new_G570 = ~new_G1238;
  assign new_G578 = ~new_G1926;
  assign new_G579 = ~new_G1921;
  assign new_G580 = ~new_G1916;
  assign new_G1256 = new_G1209 & new_G1231;
  assign new_G1261 = new_G1216 & new_G1231;
  assign new_G1266 = new_G1223 & new_G1231;
  assign new_G1271 = new_G1080 & new_G1231;
  assign new_G1486 = ~new_G1483;
  assign new_G1934 = new_G1887 & new_G1909;
  assign new_G1942 = new_G1894 & new_G1909;
  assign new_G1947 = new_G1901 & new_G1909;
  assign new_G1952 = new_G1758 & new_G1909;
  assign new_G2163 = ~new_G2160;
  assign new_G5250 = ~new_G5244;
  assign new_G3537 = ~new_G5244 | ~new_G5251;
  assign new_G5258 = ~new_G5252;
  assign new_G3542 = ~new_G5252 | ~new_G5259;
  assign new_G3782 = new_G3765 & new_G1253 & new_G3737;
  assign new_G3785 = new_G3765 & new_G1248 & new_G3737;
  assign new_G3788 = new_G3765 & new_G1243 & new_G3737;
  assign new_G3790 = new_G3780 | new_G3778 | new_G3779;
  assign new_G3843 = new_G3823 & new_G1926 & new_G3795;
  assign new_G3846 = new_G3823 & new_G1921 & new_G3795;
  assign new_G3849 = new_G3841 | new_G3839 | new_G3840;
  assign new_G3960 = ~new_G5409 | ~new_G5412;
  assign new_G5413 = ~new_G5409;
  assign new_G3963 = ~new_G5417 | ~new_G5420;
  assign new_G4010 = new_G3998 & new_G1238 & new_G3972;
  assign new_G4068 = new_G4056 & new_G1916 & new_G4030;
  assign new_G4358 = ~new_G4356 | ~new_G4357;
  assign new_G4416 = ~new_G4414 | ~new_G4415;
  assign new_G4480 = ~new_G4474;
  assign new_G4483 = ~new_G4474 | ~new_G4481;
  assign new_G4568 = ~new_G4562;
  assign new_G4571 = ~new_G4562 | ~new_G4569;
  assign new_G4822 = ~new_G4820 | ~new_G4821;
  assign new_G4880 = ~new_G4878 | ~new_G4879;
  assign new_G4938 = ~new_G4936 | ~new_G4937;
  assign new_G5022 = ~new_G5016;
  assign new_G5025 = ~new_G5016 | ~new_G5023;
  assign new_G1258 = new_G1256 | new_G1257;
  assign new_G1263 = new_G1261 | new_G1262;
  assign new_G1268 = new_G1266 | new_G1267;
  assign new_G1273 = new_G1271 | new_G1272;
  assign new_G1936 = new_G1934 | new_G1935;
  assign new_G1944 = new_G1942 | new_G1943;
  assign new_G1949 = new_G1947 | new_G1948;
  assign new_G1954 = new_G1952 | new_G1953;
  assign new_G3536 = ~new_G5247 | ~new_G5250;
  assign new_G3541 = ~new_G5255 | ~new_G5258;
  assign new_G3791 = new_G3783 | new_G3781 | new_G3782;
  assign new_G3792 = new_G3786 | new_G3784 | new_G3785;
  assign new_G3793 = new_G3789 | new_G3787 | new_G3788;
  assign new_G3850 = new_G3844 | new_G3842 | new_G3843;
  assign new_G3851 = new_G3847 | new_G3845 | new_G3846;
  assign new_G3961 = ~new_G5406 | ~new_G5413;
  assign new_G3965 = ~new_G3963 | ~new_G3964;
  assign new_G4024 = new_G4011 | new_G4009 | new_G4010;
  assign new_G4082 = new_G4069 | new_G4067 | new_G4068;
  assign new_G4482 = ~new_G4477 | ~new_G4480;
  assign new_G4570 = ~new_G4565 | ~new_G4568;
  assign new_G5024 = ~new_G5019 | ~new_G5022;
  assign new_G1666 = new_G1645 & new_G3790 & new_G1609;
  assign new_G1670 = new_G1645 & new_G3849 & new_G1621;
  assign new_G2337 = new_G2316 & new_G3790 & new_G2281;
  assign new_G2341 = new_G2316 & new_G3849 & new_G2293;
  assign new_G719 = new_G2454 & new_G3790 & new_G2418;
  assign new_G758 = new_G2454 & new_G3849 & new_G2430;
  assign new_G798 = new_G2512 & new_G3849 & new_G2488;
  assign G838 = ~new_G3849;
  assign new_G856 = new_G2512 & new_G3790 & new_G2476;
  assign G861 = ~new_G3790;
  assign new_G3538 = ~new_G3536 | ~new_G3537;
  assign new_G3543 = ~new_G3541 | ~new_G3542;
  assign new_G3962 = ~new_G3960 | ~new_G3961;
  assign new_G4364 = ~new_G4358;
  assign new_G4367 = ~new_G4358 | ~new_G4365;
  assign new_G4422 = ~new_G4416;
  assign new_G4425 = ~new_G4416 | ~new_G4423;
  assign new_G4484 = ~new_G4482 | ~new_G4483;
  assign new_G4572 = ~new_G4570 | ~new_G4571;
  assign new_G4828 = ~new_G4822;
  assign new_G4831 = ~new_G4822 | ~new_G4829;
  assign new_G4886 = ~new_G4880;
  assign new_G4889 = ~new_G4880 | ~new_G4887;
  assign new_G4944 = ~new_G4938;
  assign new_G4947 = ~new_G4938 | ~new_G4945;
  assign new_G5026 = ~new_G5024 | ~new_G5025;
  assign new_G571 = ~new_G1273;
  assign new_G572 = ~new_G1268;
  assign new_G573 = ~new_G1263;
  assign new_G574 = ~new_G1258;
  assign new_G581 = ~new_G1954;
  assign new_G582 = ~new_G1949;
  assign new_G583 = ~new_G1944;
  assign new_G584 = ~new_G1936;
  assign G623 = ~new_G1936;
  assign new_G1576 = new_G1564 & new_G4082 & new_G1540;
  assign new_G1578 = new_G1564 & new_G4024 & new_G1528;
  assign new_G659 = new_G1668 | new_G1667 | new_G1664 | new_G1666;
  assign new_G1672 = new_G1645 & new_G3791 & new_G1609;
  assign new_G1676 = new_G1645 & new_G3850 & new_G1621;
  assign new_G1678 = new_G1645 & new_G3792 & new_G1609;
  assign new_G1682 = new_G1645 & new_G3851 & new_G1621;
  assign new_G1684 = new_G1645 & new_G3793 & new_G1609;
  assign new_G2250 = new_G2238 & new_G4082 & new_G2215;
  assign new_G2252 = new_G2238 & new_G4024 & new_G2203;
  assign new_G691 = new_G2339 | new_G2338 | new_G2335 | new_G2337;
  assign new_G2343 = new_G2316 & new_G3791 & new_G2281;
  assign new_G2347 = new_G2316 & new_G3850 & new_G2293;
  assign new_G2349 = new_G2316 & new_G3792 & new_G2281;
  assign new_G2353 = new_G2316 & new_G3851 & new_G2293;
  assign new_G2355 = new_G2316 & new_G3793 & new_G2281;
  assign G722 = new_G721 | new_G720 | new_G718 | new_G719;
  assign new_G743 = new_G3594 & new_G4082 & new_G3570;
  assign new_G744 = new_G3594 & new_G4024 & new_G3558;
  assign new_G748 = new_G2454 & new_G3851 & new_G2430;
  assign new_G749 = new_G2454 & new_G3793 & new_G2418;
  assign new_G753 = new_G2454 & new_G3850 & new_G2430;
  assign new_G754 = new_G2454 & new_G3792 & new_G2418;
  assign new_G759 = new_G2454 & new_G3791 & new_G2418;
  assign new_G783 = new_G3696 & new_G4082 & new_G3672;
  assign new_G784 = new_G3696 & new_G4024 & new_G3660;
  assign new_G788 = new_G2512 & new_G3851 & new_G2488;
  assign new_G789 = new_G2512 & new_G3793 & new_G2476;
  assign new_G793 = new_G2512 & new_G3850 & new_G2488;
  assign new_G794 = new_G2512 & new_G3792 & new_G2476;
  assign new_G799 = new_G2512 & new_G3791 & new_G2476;
  assign new_G3735 = G3717 & new_G1936 & G3724;
  assign G832 = ~new_G4082;
  assign G834 = ~new_G3851;
  assign G836 = ~new_G3850;
  assign new_G3835 = ~new_G3965;
  assign G859 = new_G858 | new_G857 | new_G855 | new_G856;
  assign G871 = ~new_G4024;
  assign G873 = ~new_G3793;
  assign G875 = ~new_G3792;
  assign G877 = ~new_G3791;
  assign G998 = new_G3538;
  assign G1000 = new_G3543;
  assign new_G3651 = new_G3965 & new_G3632;
  assign new_G4013 = new_G3998 & new_G1273 & new_G3972;
  assign new_G4016 = new_G3998 & new_G1268 & new_G3972;
  assign new_G4019 = new_G3998 & new_G1263 & new_G3972;
  assign new_G4022 = new_G3998 & new_G1258 & new_G3972;
  assign new_G4071 = new_G4056 & new_G1954 & new_G4030;
  assign new_G4074 = new_G4056 & new_G1949 & new_G4030;
  assign new_G4077 = new_G4056 & new_G1944 & new_G4030;
  assign new_G4080 = new_G4056 & new_G1936 & new_G4030;
  assign new_G4096 = ~new_G4113 | ~new_G1936;
  assign new_G4366 = ~new_G4361 | ~new_G4364;
  assign new_G4424 = ~new_G4419 | ~new_G4422;
  assign new_G4830 = ~new_G4825 | ~new_G4828;
  assign new_G4888 = ~new_G4883 | ~new_G4886;
  assign new_G4946 = ~new_G4941 | ~new_G4944;
  assign G575 = new_G574 & new_G573 & new_G572 & new_G571 & new_G570 & new_G569 & new_G568 & new_G566 & new_G567;
  assign G585 = new_G584 & new_G583 & new_G582 & new_G581 & new_G580 & new_G579 & new_G578 & new_G576 & new_G577;
  assign new_G640 = new_G1580 | new_G1579 | new_G1576 | new_G1578;
  assign G661 = new_G659 & new_G1606;
  assign new_G662 = new_G1674 | new_G1673 | new_G1670 | new_G1672;
  assign new_G665 = new_G1680 | new_G1679 | new_G1676 | new_G1678;
  assign new_G668 = new_G1686 | new_G1685 | new_G1682 | new_G1684;
  assign new_G674 = new_G2254 | new_G2253 | new_G2250 | new_G2252;
  assign G693 = new_G691 & new_G2279;
  assign new_G694 = new_G2345 | new_G2344 | new_G2341 | new_G2343;
  assign new_G697 = new_G2351 | new_G2350 | new_G2347 | new_G2349;
  assign new_G700 = new_G2357 | new_G2356 | new_G2353 | new_G2355;
  assign G747 = new_G746 | new_G745 | new_G743 | new_G744;
  assign G752 = new_G751 | new_G750 | new_G748 | new_G749;
  assign G757 = new_G756 | new_G755 | new_G753 | new_G754;
  assign G762 = new_G761 | new_G760 | new_G758 | new_G759;
  assign G787 = new_G786 | new_G785 | new_G783 | new_G784;
  assign G792 = new_G791 | new_G790 | new_G788 | new_G789;
  assign G797 = new_G796 | new_G795 | new_G793 | new_G794;
  assign G802 = new_G801 | new_G800 | new_G798 | new_G799;
  assign new_G817 = new_G3735 | new_G3734 | new_G3731 | new_G3733;
  assign new_G839 = new_G3823 & new_G3835 & new_G3803;
  assign new_G3540 = ~new_G3538;
  assign new_G3545 = ~new_G3543;
  assign new_G3777 = ~new_G3962;
  assign new_G3648 = new_G3962 & new_G3632;
  assign new_G4025 = new_G4014 | new_G4012 | new_G4013;
  assign new_G4026 = new_G4017 | new_G4015 | new_G4016;
  assign new_G4027 = new_G4020 | new_G4018 | new_G4019;
  assign new_G4028 = new_G4023 | new_G4021 | new_G4022;
  assign new_G4083 = new_G4072 | new_G4070 | new_G4071;
  assign new_G4084 = new_G4075 | new_G4073 | new_G4074;
  assign new_G4085 = new_G4078 | new_G4076 | new_G4077;
  assign new_G4086 = new_G4081 | new_G4079 | new_G4080;
  assign new_G4368 = ~new_G4366 | ~new_G4367;
  assign new_G4426 = ~new_G4424 | ~new_G4425;
  assign new_G4490 = ~new_G4484;
  assign new_G4493 = ~new_G4484 | ~new_G4491;
  assign new_G4578 = ~new_G4572;
  assign new_G4581 = ~new_G4572 | ~new_G4579;
  assign new_G4832 = ~new_G4830 | ~new_G4831;
  assign new_G4890 = ~new_G4888 | ~new_G4889;
  assign new_G4948 = ~new_G4946 | ~new_G4947;
  assign new_G5032 = ~new_G5026;
  assign new_G5035 = ~new_G5026 | ~new_G5033;
  assign G642 = new_G640 & new_G1526;
  assign G664 = new_G662 & new_G1606;
  assign G667 = new_G665 & new_G1606;
  assign G670 = new_G668 & new_G1606;
  assign G676 = new_G674 & new_G2202;
  assign G696 = new_G694 & new_G2279;
  assign G699 = new_G697 & new_G2279;
  assign G702 = new_G700 & new_G2279;
  assign new_G811 = new_G4113 & new_G4096;
  assign new_G812 = new_G4096 & new_G1936;
  assign G818 = new_G816 & new_G817;
  assign new_G853 = new_G3970 & new_G3535 & new_G3545 & G562 & new_G3540;
  assign new_G878 = new_G3765 & new_G3777 & new_G3745;
  assign new_G4492 = ~new_G4487 | ~new_G4490;
  assign new_G4580 = ~new_G4575 | ~new_G4578;
  assign new_G5034 = ~new_G5029 | ~new_G5032;
  assign new_G1582 = new_G1564 & new_G4083 & new_G1540;
  assign new_G1584 = new_G1564 & new_G4025 & new_G1528;
  assign new_G1588 = new_G1564 & new_G4084 & new_G1540;
  assign new_G1590 = new_G1564 & new_G4026 & new_G1528;
  assign new_G1594 = new_G1564 & new_G4085 & new_G1540;
  assign new_G1596 = new_G1564 & new_G4027 & new_G1528;
  assign new_G1600 = new_G1564 & new_G4086 & new_G1540;
  assign new_G1602 = new_G1564 & new_G4028 & new_G1528;
  assign new_G2256 = new_G2238 & new_G4083 & new_G2215;
  assign new_G2258 = new_G2238 & new_G4025 & new_G2203;
  assign new_G2262 = new_G2238 & new_G4084 & new_G2215;
  assign new_G2264 = new_G2238 & new_G4026 & new_G2203;
  assign new_G2268 = new_G2238 & new_G4085 & new_G2215;
  assign new_G2270 = new_G2238 & new_G4027 & new_G2203;
  assign new_G2274 = new_G2238 & new_G4086 & new_G2215;
  assign new_G2276 = new_G2238 & new_G4028 & new_G2203;
  assign new_G708 = new_G3696 & new_G4086 & new_G3672;
  assign new_G709 = new_G3696 & new_G4028 & new_G3660;
  assign new_G723 = new_G3594 & new_G4086 & new_G3570;
  assign new_G724 = new_G3594 & new_G4028 & new_G3558;
  assign new_G728 = new_G3594 & new_G4085 & new_G3570;
  assign new_G729 = new_G3594 & new_G4027 & new_G3558;
  assign new_G733 = new_G3594 & new_G4084 & new_G3570;
  assign new_G734 = new_G3594 & new_G4026 & new_G3558;
  assign new_G738 = new_G3594 & new_G4083 & new_G3570;
  assign new_G739 = new_G3594 & new_G4025 & new_G3558;
  assign new_G768 = new_G3696 & new_G4085 & new_G3672;
  assign new_G769 = new_G3696 & new_G4027 & new_G3660;
  assign new_G773 = new_G3696 & new_G4084 & new_G3672;
  assign new_G774 = new_G3696 & new_G4026 & new_G3660;
  assign new_G778 = new_G3696 & new_G4083 & new_G3672;
  assign new_G779 = new_G3696 & new_G4025 & new_G3660;
  assign G813 = new_G811 | new_G812;
  assign G824 = ~new_G4086;
  assign G826 = ~new_G4085;
  assign G828 = ~new_G4084;
  assign G830 = ~new_G4083;
  assign G854 = G245 & new_G852 & new_G853;
  assign G863 = ~new_G4028;
  assign G865 = ~new_G4027;
  assign G867 = ~new_G4026;
  assign G869 = ~new_G4025;
  assign new_G4374 = ~new_G4368;
  assign new_G4377 = ~new_G4368 | ~new_G4375;
  assign new_G4432 = ~new_G4426;
  assign new_G4435 = ~new_G4426 | ~new_G4433;
  assign new_G4494 = ~new_G4492 | ~new_G4493;
  assign new_G4582 = ~new_G4580 | ~new_G4581;
  assign new_G4838 = ~new_G4832;
  assign new_G4841 = ~new_G4832 | ~new_G4839;
  assign new_G4896 = ~new_G4890;
  assign new_G4899 = ~new_G4890 | ~new_G4897;
  assign new_G4954 = ~new_G4948;
  assign new_G4957 = ~new_G4948 | ~new_G4955;
  assign new_G5036 = ~new_G5034 | ~new_G5035;
  assign new_G643 = new_G1586 | new_G1585 | new_G1582 | new_G1584;
  assign new_G646 = new_G1592 | new_G1591 | new_G1588 | new_G1590;
  assign new_G649 = new_G1598 | new_G1597 | new_G1594 | new_G1596;
  assign new_G652 = new_G1604 | new_G1603 | new_G1600 | new_G1602;
  assign new_G677 = new_G2260 | new_G2259 | new_G2256 | new_G2258;
  assign new_G680 = new_G2266 | new_G2265 | new_G2262 | new_G2264;
  assign new_G683 = new_G2272 | new_G2271 | new_G2268 | new_G2270;
  assign new_G686 = new_G2278 | new_G2277 | new_G2274 | new_G2276;
  assign G712 = new_G711 | new_G710 | new_G708 | new_G709;
  assign G727 = new_G726 | new_G725 | new_G723 | new_G724;
  assign G732 = new_G731 | new_G730 | new_G728 | new_G729;
  assign G737 = new_G736 | new_G735 | new_G733 | new_G734;
  assign G742 = new_G741 | new_G740 | new_G738 | new_G739;
  assign G772 = new_G771 | new_G770 | new_G768 | new_G769;
  assign G777 = new_G776 | new_G775 | new_G773 | new_G774;
  assign G782 = new_G781 | new_G780 | new_G778 | new_G779;
  assign new_G4376 = ~new_G4371 | ~new_G4374;
  assign new_G4434 = ~new_G4429 | ~new_G4432;
  assign new_G4840 = ~new_G4835 | ~new_G4838;
  assign new_G4898 = ~new_G4893 | ~new_G4896;
  assign new_G4956 = ~new_G4951 | ~new_G4954;
  assign G645 = new_G643 & new_G1526;
  assign G648 = new_G646 & new_G1526;
  assign G651 = new_G649 & new_G1526;
  assign G654 = new_G652 & new_G1526;
  assign G679 = new_G677 & new_G2202;
  assign G682 = new_G680 & new_G2202;
  assign G685 = new_G683 & new_G2202;
  assign G688 = new_G686 & new_G2202;
  assign new_G4378 = ~new_G4376 | ~new_G4377;
  assign new_G4436 = ~new_G4434 | ~new_G4435;
  assign new_G4500 = ~new_G4494;
  assign new_G4503 = ~new_G4494 | ~new_G4501;
  assign new_G4588 = ~new_G4582;
  assign new_G4591 = ~new_G4582 | ~new_G4589;
  assign new_G4842 = ~new_G4840 | ~new_G4841;
  assign new_G4900 = ~new_G4898 | ~new_G4899;
  assign new_G4958 = ~new_G4956 | ~new_G4957;
  assign new_G5042 = ~new_G5036;
  assign new_G5045 = ~new_G5036 | ~new_G5043;
  assign new_G4502 = ~new_G4497 | ~new_G4500;
  assign new_G4590 = ~new_G4585 | ~new_G4588;
  assign new_G5044 = ~new_G5039 | ~new_G5042;
  assign new_G4384 = ~new_G4378;
  assign new_G4387 = ~new_G4378 | ~new_G4385;
  assign new_G4442 = ~new_G4436;
  assign new_G4445 = ~new_G4436 | ~new_G4443;
  assign new_G4504 = ~new_G4502 | ~new_G4503;
  assign new_G4592 = ~new_G4590 | ~new_G4591;
  assign new_G4848 = ~new_G4842;
  assign new_G4851 = ~new_G4842 | ~new_G4849;
  assign new_G4906 = ~new_G4900;
  assign new_G4909 = ~new_G4900 | ~new_G4907;
  assign new_G4964 = ~new_G4958;
  assign new_G4967 = ~new_G4958 | ~new_G4965;
  assign new_G5046 = ~new_G5044 | ~new_G5045;
  assign new_G4386 = ~new_G4381 | ~new_G4384;
  assign new_G4444 = ~new_G4439 | ~new_G4442;
  assign new_G4850 = ~new_G4845 | ~new_G4848;
  assign new_G4908 = ~new_G4903 | ~new_G4906;
  assign new_G4966 = ~new_G4961 | ~new_G4964;
  assign new_G4388 = ~new_G4386 | ~new_G4387;
  assign new_G4446 = ~new_G4444 | ~new_G4445;
  assign new_G4510 = ~new_G4504;
  assign new_G4513 = ~new_G4504 | ~new_G4511;
  assign new_G4598 = ~new_G4592;
  assign new_G4601 = ~new_G4592 | ~new_G4599;
  assign new_G4852 = ~new_G4850 | ~new_G4851;
  assign new_G4910 = ~new_G4908 | ~new_G4909;
  assign new_G4968 = ~new_G4966 | ~new_G4967;
  assign new_G5052 = ~new_G5046;
  assign new_G5055 = ~new_G5046 | ~new_G5053;
  assign new_G4512 = ~new_G4507 | ~new_G4510;
  assign new_G4600 = ~new_G4595 | ~new_G4598;
  assign new_G5054 = ~new_G5049 | ~new_G5052;
  assign new_G4394 = ~new_G4388;
  assign new_G4397 = ~new_G4388 | ~new_G4395;
  assign new_G4452 = ~new_G4446;
  assign new_G4455 = ~new_G4446 | ~new_G4453;
  assign new_G4514 = ~new_G4512 | ~new_G4513;
  assign new_G4602 = ~new_G4600 | ~new_G4601;
  assign new_G4858 = ~new_G4852;
  assign new_G4861 = ~new_G4852 | ~new_G4859;
  assign new_G4916 = ~new_G4910;
  assign new_G4919 = ~new_G4910 | ~new_G4917;
  assign new_G4974 = ~new_G4968;
  assign new_G4977 = ~new_G4968 | ~new_G4975;
  assign new_G5056 = ~new_G5054 | ~new_G5055;
  assign new_G4396 = ~new_G4391 | ~new_G4394;
  assign new_G4454 = ~new_G4449 | ~new_G4452;
  assign new_G4860 = ~new_G4855 | ~new_G4858;
  assign new_G4918 = ~new_G4913 | ~new_G4916;
  assign new_G4976 = ~new_G4971 | ~new_G4974;
  assign new_G4398 = ~new_G4396 | ~new_G4397;
  assign new_G4456 = ~new_G4454 | ~new_G4455;
  assign new_G4520 = ~new_G4514;
  assign new_G4523 = ~new_G4514 | ~new_G4521;
  assign new_G4608 = ~new_G4602;
  assign new_G4611 = ~new_G4602 | ~new_G4609;
  assign new_G4862 = ~new_G4860 | ~new_G4861;
  assign new_G4920 = ~new_G4918 | ~new_G4919;
  assign new_G4978 = ~new_G4976 | ~new_G4977;
  assign new_G5062 = ~new_G5056;
  assign new_G5065 = ~new_G5056 | ~new_G5063;
  assign new_G4522 = ~new_G4517 | ~new_G4520;
  assign new_G4610 = ~new_G4605 | ~new_G4608;
  assign new_G5064 = ~new_G5059 | ~new_G5062;
  assign new_G4404 = ~new_G4398;
  assign new_G1488 = ~new_G4398 | ~new_G4405;
  assign new_G4462 = ~new_G4456;
  assign new_G1493 = ~new_G4456 | ~new_G4463;
  assign new_G4868 = ~new_G4862;
  assign new_G2165 = ~new_G4862 | ~new_G4869;
  assign new_G4926 = ~new_G4920;
  assign new_G2170 = ~new_G4920 | ~new_G4927;
  assign new_G4524 = ~new_G4522 | ~new_G4523;
  assign new_G4612 = ~new_G4610 | ~new_G4611;
  assign new_G4984 = ~new_G4978;
  assign new_G4987 = ~new_G4978 | ~new_G4985;
  assign new_G5066 = ~new_G5064 | ~new_G5065;
  assign new_G1487 = ~new_G4401 | ~new_G4404;
  assign new_G1492 = ~new_G4459 | ~new_G4462;
  assign new_G2164 = ~new_G4865 | ~new_G4868;
  assign new_G2169 = ~new_G4923 | ~new_G4926;
  assign new_G4986 = ~new_G4981 | ~new_G4984;
  assign new_G1489 = ~new_G1487 | ~new_G1488;
  assign new_G1494 = ~new_G1492 | ~new_G1493;
  assign new_G2166 = ~new_G2164 | ~new_G2165;
  assign new_G2171 = ~new_G2169 | ~new_G2170;
  assign new_G4530 = ~new_G4524;
  assign new_G4533 = ~new_G4524 | ~new_G4531;
  assign new_G4618 = ~new_G4612;
  assign new_G4543 = ~new_G4612 | ~new_G4619;
  assign new_G4988 = ~new_G4986 | ~new_G4987;
  assign new_G5072 = ~new_G5066;
  assign new_G4997 = ~new_G5066 | ~new_G5073;
  assign new_G4532 = ~new_G4527 | ~new_G4530;
  assign new_G4542 = ~new_G4615 | ~new_G4618;
  assign new_G4996 = ~new_G5069 | ~new_G5072;
  assign new_G1513 = new_G1502 & new_G1494 & new_G1462;
  assign new_G1514 = new_G1502 & new_G1489 & new_G1458;
  assign new_G1515 = G1497 & new_G1494 & new_G1483;
  assign new_G1516 = G1497 & new_G1489 & new_G1486;
  assign new_G4994 = ~new_G4988;
  assign new_G2184 = ~new_G4988 | ~new_G4995;
  assign new_G2190 = new_G2179 & new_G2171 & new_G2139;
  assign new_G2191 = new_G2179 & new_G2166 & new_G2135;
  assign new_G2192 = G2174 & new_G2171 & new_G2160;
  assign new_G2193 = G2174 & new_G2166 & new_G2163;
  assign new_G4534 = ~new_G4532 | ~new_G4533;
  assign new_G4544 = ~new_G4542 | ~new_G4543;
  assign new_G4998 = ~new_G4996 | ~new_G4997;
  assign new_G2183 = ~new_G4991 | ~new_G4994;
  assign new_G4620 = new_G1516 | new_G1515 | new_G1513 | new_G1514;
  assign new_G5074 = new_G2193 | new_G2192 | new_G2190 | new_G2191;
  assign new_G4540 = ~new_G4534;
  assign new_G1507 = ~new_G4534 | ~new_G4541;
  assign new_G4550 = ~new_G4544;
  assign new_G1510 = ~new_G4544 | ~new_G4551;
  assign new_G2185 = ~new_G2183 | ~new_G2184;
  assign new_G5004 = ~new_G4998;
  assign new_G2187 = ~new_G4998 | ~new_G5005;
  assign new_G1506 = ~new_G4537 | ~new_G4540;
  assign new_G1509 = ~new_G4547 | ~new_G4550;
  assign new_G4626 = ~new_G4620;
  assign new_G2186 = ~new_G5001 | ~new_G5004;
  assign new_G2195 = G2174 & new_G2185;
  assign new_G5080 = ~new_G5074;
  assign new_G1508 = ~new_G1506 | ~new_G1507;
  assign new_G1511 = ~new_G1509 | ~new_G1510;
  assign new_G2188 = ~new_G2186 | ~new_G2187;
  assign new_G1512 = ~new_G1511;
  assign new_G1518 = G1497 & new_G1508;
  assign new_G2189 = ~new_G2188;
  assign new_G1517 = new_G1512 & new_G1502;
  assign new_G2194 = new_G2189 & new_G2179;
  assign new_G4623 = new_G1517 | new_G1518;
  assign new_G5077 = new_G2194 | new_G2195;
  assign new_G1519 = ~new_G4623 | ~new_G4626;
  assign new_G4627 = ~new_G4623;
  assign new_G2196 = ~new_G5077 | ~new_G5080;
  assign new_G5081 = ~new_G5077;
  assign new_G1520 = ~new_G4620 | ~new_G4627;
  assign new_G2197 = ~new_G5074 | ~new_G5081;
  assign new_G1521 = ~new_G1519 | ~new_G1520;
  assign new_G2198 = ~new_G2196 | ~new_G2197;
  assign new_G840 = new_G3823 & new_G2198 & new_G3795;
  assign new_G879 = new_G3765 & new_G1521 & new_G3737;
  assign new_G1524 = ~new_G1521;
  assign new_G2201 = ~new_G2198;
  assign G843 = new_G842 | new_G841 | new_G839 | new_G840;
  assign G882 = new_G881 | new_G880 | new_G878 | new_G879;
  assign new_G3649 = new_G1524 & new_G3628;
  assign new_G3652 = new_G2201 & new_G3628;
  assign new_G3657 = new_G3648 | new_G3649;
  assign new_G3658 = new_G3651 | new_G3652;
  assign new_G3636 = new_G3657 & new_G3622;
  assign new_G3639 = new_G3658 & new_G3622;
  assign new_G3642 = new_G3657 & new_G3622;
  assign new_G3645 = new_G3658 & new_G3622;
  assign new_G3653 = new_G3636 | new_G3637;
  assign new_G3654 = new_G3639 | new_G3640;
  assign new_G3655 = new_G3642 | new_G3643;
  assign new_G3656 = new_G3645 | new_G3646;
  assign new_G763 = new_G2454 & new_G3656 & new_G2430;
  assign new_G764 = new_G2454 & new_G3655 & new_G2418;
  assign new_G803 = new_G2512 & new_G3656 & new_G2488;
  assign new_G804 = new_G2512 & new_G3655 & new_G2476;
  assign new_G1657 = new_G1645 & new_G3654 & new_G1621;
  assign new_G1659 = new_G1645 & new_G3653 & new_G1609;
  assign new_G2328 = new_G2316 & new_G3654 & new_G2293;
  assign new_G2330 = new_G2316 & new_G3653 & new_G2281;
  assign new_G1662 = new_G1661 | new_G1660 | new_G1657 | new_G1659;
  assign new_G2333 = new_G2332 | new_G2331 | new_G2328 | new_G2330;
  assign G767 = new_G766 | new_G765 | new_G763 | new_G764;
  assign G807 = new_G806 | new_G805 | new_G803 | new_G804;
  assign new_G657 = new_G1662 & new_G1606;
  assign new_G689 = new_G2333 & new_G2279;
  assign G658 = ~new_G657;
  assign G690 = ~new_G689;
endmodule
