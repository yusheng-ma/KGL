// Benchmark "./benchmarks/iscas85/c6288" written by ABC on Sun Apr 28 12:32:39 2024

module c6288  ( 
    G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire new_G546gat, new_G549gat, new_G552gat, new_G555gat, new_G558gat,
    new_G561gat, new_G564gat, new_G567gat, new_G570gat, new_G573gat,
    new_G576gat, new_G579gat, new_G582gat, new_G585gat, new_G588gat,
    new_G591gat, new_G594gat, new_G597gat, new_G600gat, new_G603gat,
    new_G606gat, new_G609gat, new_G612gat, new_G615gat, new_G618gat,
    new_G621gat, new_G624gat, new_G627gat, new_G630gat, new_G633gat,
    new_G636gat, new_G639gat, new_G642gat, new_G645gat, new_G648gat,
    new_G651gat, new_G654gat, new_G657gat, new_G660gat, new_G663gat,
    new_G666gat, new_G669gat, new_G672gat, new_G675gat, new_G678gat,
    new_G681gat, new_G684gat, new_G687gat, new_G690gat, new_G693gat,
    new_G696gat, new_G699gat, new_G702gat, new_G705gat, new_G708gat,
    new_G711gat, new_G714gat, new_G717gat, new_G720gat, new_G723gat,
    new_G726gat, new_G729gat, new_G732gat, new_G735gat, new_G738gat,
    new_G741gat, new_G744gat, new_G747gat, new_G750gat, new_G753gat,
    new_G756gat, new_G759gat, new_G762gat, new_G765gat, new_G768gat,
    new_G771gat, new_G774gat, new_G777gat, new_G780gat, new_G783gat,
    new_G786gat, new_G789gat, new_G792gat, new_G795gat, new_G798gat,
    new_G801gat, new_G804gat, new_G807gat, new_G810gat, new_G813gat,
    new_G816gat, new_G819gat, new_G822gat, new_G825gat, new_G828gat,
    new_G831gat, new_G834gat, new_G837gat, new_G840gat, new_G843gat,
    new_G846gat, new_G849gat, new_G852gat, new_G855gat, new_G858gat,
    new_G861gat, new_G864gat, new_G867gat, new_G870gat, new_G873gat,
    new_G876gat, new_G879gat, new_G882gat, new_G885gat, new_G888gat,
    new_G891gat, new_G894gat, new_G897gat, new_G900gat, new_G903gat,
    new_G906gat, new_G909gat, new_G912gat, new_G915gat, new_G918gat,
    new_G921gat, new_G924gat, new_G927gat, new_G930gat, new_G933gat,
    new_G936gat, new_G939gat, new_G942gat, new_G945gat, new_G948gat,
    new_G951gat, new_G954gat, new_G957gat, new_G960gat, new_G963gat,
    new_G966gat, new_G969gat, new_G972gat, new_G975gat, new_G978gat,
    new_G981gat, new_G984gat, new_G987gat, new_G990gat, new_G993gat,
    new_G996gat, new_G999gat, new_G1002gat, new_G1005gat, new_G1008gat,
    new_G1011gat, new_G1014gat, new_G1017gat, new_G1020gat, new_G1023gat,
    new_G1026gat, new_G1029gat, new_G1032gat, new_G1035gat, new_G1038gat,
    new_G1041gat, new_G1044gat, new_G1047gat, new_G1050gat, new_G1053gat,
    new_G1056gat, new_G1059gat, new_G1062gat, new_G1065gat, new_G1068gat,
    new_G1071gat, new_G1074gat, new_G1077gat, new_G1080gat, new_G1083gat,
    new_G1086gat, new_G1089gat, new_G1092gat, new_G1095gat, new_G1098gat,
    new_G1101gat, new_G1104gat, new_G1107gat, new_G1110gat, new_G1113gat,
    new_G1116gat, new_G1119gat, new_G1122gat, new_G1125gat, new_G1128gat,
    new_G1131gat, new_G1134gat, new_G1137gat, new_G1140gat, new_G1143gat,
    new_G1146gat, new_G1149gat, new_G1152gat, new_G1155gat, new_G1158gat,
    new_G1161gat, new_G1164gat, new_G1167gat, new_G1170gat, new_G1173gat,
    new_G1176gat, new_G1179gat, new_G1182gat, new_G1185gat, new_G1188gat,
    new_G1191gat, new_G1194gat, new_G1197gat, new_G1200gat, new_G1203gat,
    new_G1206gat, new_G1209gat, new_G1212gat, new_G1215gat, new_G1218gat,
    new_G1221gat, new_G1224gat, new_G1227gat, new_G1230gat, new_G1233gat,
    new_G1236gat, new_G1239gat, new_G1242gat, new_G1245gat, new_G1248gat,
    new_G1251gat, new_G1254gat, new_G1257gat, new_G1260gat, new_G1263gat,
    new_G1266gat, new_G1269gat, new_G1272gat, new_G1275gat, new_G1278gat,
    new_G1281gat, new_G1284gat, new_G1287gat, new_G1290gat, new_G1293gat,
    new_G1296gat, new_G1299gat, new_G1302gat, new_G1305gat, new_G1308gat,
    new_G1311gat, new_G1315gat, new_G1319gat, new_G1323gat, new_G1327gat,
    new_G1331gat, new_G1335gat, new_G1339gat, new_G1343gat, new_G1347gat,
    new_G1351gat, new_G1355gat, new_G1359gat, new_G1363gat, new_G1367gat,
    new_G1371gat, new_G1372gat, new_G1373gat, new_G1374gat, new_G1375gat,
    new_G1376gat, new_G1377gat, new_G1378gat, new_G1379gat, new_G1380gat,
    new_G1381gat, new_G1382gat, new_G1383gat, new_G1384gat, new_G1385gat,
    new_G1386gat, new_G1387gat, new_G1388gat, new_G1389gat, new_G1390gat,
    new_G1391gat, new_G1392gat, new_G1393gat, new_G1394gat, new_G1395gat,
    new_G1396gat, new_G1397gat, new_G1398gat, new_G1399gat, new_G1400gat,
    new_G1401gat, new_G1404gat, new_G1407gat, new_G1410gat, new_G1413gat,
    new_G1416gat, new_G1419gat, new_G1422gat, new_G1425gat, new_G1428gat,
    new_G1431gat, new_G1434gat, new_G1437gat, new_G1440gat, new_G1443gat,
    new_G1446gat, new_G1450gat, new_G1454gat, new_G1458gat, new_G1462gat,
    new_G1466gat, new_G1470gat, new_G1474gat, new_G1478gat, new_G1482gat,
    new_G1486gat, new_G1490gat, new_G1494gat, new_G1498gat, new_G1502gat,
    new_G1506gat, new_G1507gat, new_G1508gat, new_G1511gat, new_G1512gat,
    new_G1513gat, new_G1516gat, new_G1517gat, new_G1518gat, new_G1521gat,
    new_G1522gat, new_G1523gat, new_G1526gat, new_G1527gat, new_G1528gat,
    new_G1531gat, new_G1532gat, new_G1533gat, new_G1536gat, new_G1537gat,
    new_G1538gat, new_G1541gat, new_G1542gat, new_G1543gat, new_G1546gat,
    new_G1547gat, new_G1548gat, new_G1551gat, new_G1552gat, new_G1553gat,
    new_G1556gat, new_G1557gat, new_G1558gat, new_G1561gat, new_G1562gat,
    new_G1563gat, new_G1566gat, new_G1567gat, new_G1568gat, new_G1571gat,
    new_G1572gat, new_G1573gat, new_G1576gat, new_G1577gat, new_G1578gat,
    new_G1582gat, new_G1585gat, new_G1588gat, new_G1591gat, new_G1594gat,
    new_G1597gat, new_G1600gat, new_G1603gat, new_G1606gat, new_G1609gat,
    new_G1612gat, new_G1615gat, new_G1618gat, new_G1621gat, new_G1624gat,
    new_G1628gat, new_G1632gat, new_G1636gat, new_G1640gat, new_G1644gat,
    new_G1648gat, new_G1652gat, new_G1656gat, new_G1660gat, new_G1664gat,
    new_G1668gat, new_G1672gat, new_G1676gat, new_G1680gat, new_G1684gat,
    new_G1685gat, new_G1686gat, new_G1687gat, new_G1688gat, new_G1689gat,
    new_G1690gat, new_G1691gat, new_G1692gat, new_G1693gat, new_G1694gat,
    new_G1695gat, new_G1696gat, new_G1697gat, new_G1698gat, new_G1699gat,
    new_G1700gat, new_G1701gat, new_G1702gat, new_G1703gat, new_G1704gat,
    new_G1705gat, new_G1706gat, new_G1707gat, new_G1708gat, new_G1709gat,
    new_G1710gat, new_G1711gat, new_G1712gat, new_G1713gat, new_G1714gat,
    new_G1717gat, new_G1720gat, new_G1723gat, new_G1726gat, new_G1729gat,
    new_G1732gat, new_G1735gat, new_G1738gat, new_G1741gat, new_G1744gat,
    new_G1747gat, new_G1750gat, new_G1753gat, new_G1756gat, new_G1759gat,
    new_G1763gat, new_G1767gat, new_G1771gat, new_G1775gat, new_G1779gat,
    new_G1783gat, new_G1787gat, new_G1791gat, new_G1795gat, new_G1799gat,
    new_G1803gat, new_G1807gat, new_G1811gat, new_G1815gat, new_G1819gat,
    new_G1820gat, new_G1821gat, new_G1824gat, new_G1825gat, new_G1826gat,
    new_G1829gat, new_G1830gat, new_G1831gat, new_G1834gat, new_G1835gat,
    new_G1836gat, new_G1839gat, new_G1840gat, new_G1841gat, new_G1844gat,
    new_G1845gat, new_G1846gat, new_G1849gat, new_G1850gat, new_G1851gat,
    new_G1854gat, new_G1855gat, new_G1856gat, new_G1859gat, new_G1860gat,
    new_G1861gat, new_G1864gat, new_G1865gat, new_G1866gat, new_G1869gat,
    new_G1870gat, new_G1871gat, new_G1874gat, new_G1875gat, new_G1876gat,
    new_G1879gat, new_G1880gat, new_G1881gat, new_G1884gat, new_G1885gat,
    new_G1886gat, new_G1889gat, new_G1890gat, new_G1891gat, new_G1894gat,
    new_G1897gat, new_G1902gat, new_G1905gat, new_G1908gat, new_G1911gat,
    new_G1914gat, new_G1917gat, new_G1920gat, new_G1923gat, new_G1926gat,
    new_G1929gat, new_G1932gat, new_G1935gat, new_G1938gat, new_G1941gat,
    new_G1945gat, new_G1946gat, new_G1947gat, new_G1951gat, new_G1955gat,
    new_G1959gat, new_G1963gat, new_G1967gat, new_G1971gat, new_G1975gat,
    new_G1979gat, new_G1983gat, new_G1987gat, new_G1991gat, new_G1995gat,
    new_G1999gat, new_G2000gat, new_G2001gat, new_G2004gat, new_G2005gat,
    new_G2006gat, new_G2007gat, new_G2008gat, new_G2009gat, new_G2010gat,
    new_G2011gat, new_G2012gat, new_G2013gat, new_G2014gat, new_G2015gat,
    new_G2016gat, new_G2017gat, new_G2018gat, new_G2019gat, new_G2020gat,
    new_G2021gat, new_G2022gat, new_G2023gat, new_G2024gat, new_G2025gat,
    new_G2026gat, new_G2027gat, new_G2028gat, new_G2029gat, new_G2030gat,
    new_G2033gat, new_G2037gat, new_G2040gat, new_G2043gat, new_G2046gat,
    new_G2049gat, new_G2052gat, new_G2055gat, new_G2058gat, new_G2061gat,
    new_G2064gat, new_G2067gat, new_G2070gat, new_G2073gat, new_G2076gat,
    new_G2080gat, new_G2081gat, new_G2082gat, new_G2085gat, new_G2089gat,
    new_G2093gat, new_G2097gat, new_G2101gat, new_G2105gat, new_G2109gat,
    new_G2113gat, new_G2117gat, new_G2121gat, new_G2125gat, new_G2129gat,
    new_G2133gat, new_G2137gat, new_G2138gat, new_G2139gat, new_G2142gat,
    new_G2145gat, new_G2149gat, new_G2150gat, new_G2151gat, new_G2154gat,
    new_G2155gat, new_G2156gat, new_G2159gat, new_G2160gat, new_G2161gat,
    new_G2164gat, new_G2165gat, new_G2166gat, new_G2169gat, new_G2170gat,
    new_G2171gat, new_G2174gat, new_G2175gat, new_G2176gat, new_G2179gat,
    new_G2180gat, new_G2181gat, new_G2184gat, new_G2185gat, new_G2186gat,
    new_G2189gat, new_G2190gat, new_G2191gat, new_G2194gat, new_G2195gat,
    new_G2196gat, new_G2199gat, new_G2200gat, new_G2201gat, new_G2204gat,
    new_G2205gat, new_G2206gat, new_G2209gat, new_G2210gat, new_G2211gat,
    new_G2214gat, new_G2217gat, new_G2221gat, new_G2222gat, new_G2224gat,
    new_G2227gat, new_G2230gat, new_G2233gat, new_G2236gat, new_G2239gat,
    new_G2242gat, new_G2245gat, new_G2248gat, new_G2251gat, new_G2254gat,
    new_G2257gat, new_G2260gat, new_G2264gat, new_G2265gat, new_G2266gat,
    new_G2269gat, new_G2273gat, new_G2277gat, new_G2281gat, new_G2285gat,
    new_G2289gat, new_G2293gat, new_G2297gat, new_G2301gat, new_G2305gat,
    new_G2309gat, new_G2313gat, new_G2317gat, new_G2318gat, new_G2319gat,
    new_G2322gat, new_G2326gat, new_G2327gat, new_G2328gat, new_G2329gat,
    new_G2330gat, new_G2331gat, new_G2332gat, new_G2333gat, new_G2334gat,
    new_G2335gat, new_G2336gat, new_G2337gat, new_G2338gat, new_G2339gat,
    new_G2340gat, new_G2341gat, new_G2342gat, new_G2343gat, new_G2344gat,
    new_G2345gat, new_G2346gat, new_G2347gat, new_G2348gat, new_G2349gat,
    new_G2350gat, new_G2353gat, new_G2357gat, new_G2358gat, new_G2359gat,
    new_G2362gat, new_G2365gat, new_G2368gat, new_G2371gat, new_G2374gat,
    new_G2377gat, new_G2380gat, new_G2383gat, new_G2386gat, new_G2389gat,
    new_G2392gat, new_G2395gat, new_G2398gat, new_G2402gat, new_G2403gat,
    new_G2404gat, new_G2407gat, new_G2410gat, new_G2414gat, new_G2418gat,
    new_G2422gat, new_G2426gat, new_G2430gat, new_G2434gat, new_G2438gat,
    new_G2442gat, new_G2446gat, new_G2450gat, new_G2454gat, new_G2458gat,
    new_G2462gat, new_G2463gat, new_G2464gat, new_G2467gat, new_G2470gat,
    new_G2474gat, new_G2475gat, new_G2476gat, new_G2477gat, new_G2478gat,
    new_G2481gat, new_G2482gat, new_G2483gat, new_G2486gat, new_G2487gat,
    new_G2488gat, new_G2491gat, new_G2492gat, new_G2493gat, new_G2496gat,
    new_G2497gat, new_G2498gat, new_G2501gat, new_G2502gat, new_G2503gat,
    new_G2506gat, new_G2507gat, new_G2508gat, new_G2511gat, new_G2512gat,
    new_G2513gat, new_G2516gat, new_G2517gat, new_G2518gat, new_G2521gat,
    new_G2522gat, new_G2523gat, new_G2526gat, new_G2527gat, new_G2528gat,
    new_G2531gat, new_G2532gat, new_G2533gat, new_G2536gat, new_G2539gat,
    new_G2543gat, new_G2544gat, new_G2545gat, new_G2549gat, new_G2552gat,
    new_G2555gat, new_G2558gat, new_G2561gat, new_G2564gat, new_G2567gat,
    new_G2570gat, new_G2573gat, new_G2576gat, new_G2579gat, new_G2582gat,
    new_G2586gat, new_G2587gat, new_G2588gat, new_G2591gat, new_G2595gat,
    new_G2599gat, new_G2603gat, new_G2607gat, new_G2611gat, new_G2615gat,
    new_G2619gat, new_G2623gat, new_G2627gat, new_G2631gat, new_G2635gat,
    new_G2639gat, new_G2640gat, new_G2641gat, new_G2644gat, new_G2648gat,
    new_G2649gat, new_G2650gat, new_G2653gat, new_G2654gat, new_G2655gat,
    new_G2656gat, new_G2657gat, new_G2658gat, new_G2659gat, new_G2660gat,
    new_G2661gat, new_G2662gat, new_G2663gat, new_G2664gat, new_G2665gat,
    new_G2666gat, new_G2667gat, new_G2668gat, new_G2669gat, new_G2670gat,
    new_G2671gat, new_G2672gat, new_G2673gat, new_G2674gat, new_G2675gat,
    new_G2678gat, new_G2682gat, new_G2683gat, new_G2684gat, new_G2687gat,
    new_G2690gat, new_G2694gat, new_G2697gat, new_G2700gat, new_G2703gat,
    new_G2706gat, new_G2709gat, new_G2712gat, new_G2715gat, new_G2718gat,
    new_G2721gat, new_G2724gat, new_G2727gat, new_G2731gat, new_G2732gat,
    new_G2733gat, new_G2736gat, new_G2739gat, new_G2743gat, new_G2744gat,
    new_G2745gat, new_G2749gat, new_G2753gat, new_G2757gat, new_G2761gat,
    new_G2765gat, new_G2769gat, new_G2773gat, new_G2777gat, new_G2781gat,
    new_G2785gat, new_G2789gat, new_G2790gat, new_G2791gat, new_G2794gat,
    new_G2797gat, new_G2801gat, new_G2802gat, new_G2803gat, new_G2806gat,
    new_G2807gat, new_G2808gat, new_G2811gat, new_G2812gat, new_G2813gat,
    new_G2816gat, new_G2817gat, new_G2818gat, new_G2821gat, new_G2822gat,
    new_G2823gat, new_G2826gat, new_G2827gat, new_G2828gat, new_G2831gat,
    new_G2832gat, new_G2833gat, new_G2836gat, new_G2837gat, new_G2838gat,
    new_G2841gat, new_G2842gat, new_G2843gat, new_G2846gat, new_G2847gat,
    new_G2848gat, new_G2851gat, new_G2852gat, new_G2853gat, new_G2856gat,
    new_G2857gat, new_G2858gat, new_G2861gat, new_G2864gat, new_G2868gat,
    new_G2869gat, new_G2870gat, new_G2873gat, new_G2878gat, new_G2881gat,
    new_G2884gat, new_G2887gat, new_G2890gat, new_G2893gat, new_G2896gat,
    new_G2899gat, new_G2902gat, new_G2905gat, new_G2908gat, new_G2912gat,
    new_G2913gat, new_G2914gat, new_G2917gat, new_G2921gat, new_G2922gat,
    new_G2923gat, new_G2926gat, new_G2930gat, new_G2934gat, new_G2938gat,
    new_G2942gat, new_G2946gat, new_G2950gat, new_G2954gat, new_G2958gat,
    new_G2962gat, new_G2966gat, new_G2967gat, new_G2968gat, new_G2971gat,
    new_G2975gat, new_G2976gat, new_G2977gat, new_G2980gat, new_G2983gat,
    new_G2987gat, new_G2988gat, new_G2989gat, new_G2990gat, new_G2991gat,
    new_G2992gat, new_G2993gat, new_G2994gat, new_G2995gat, new_G2996gat,
    new_G2997gat, new_G2998gat, new_G2999gat, new_G3000gat, new_G3001gat,
    new_G3002gat, new_G3003gat, new_G3004gat, new_G3005gat, new_G3006gat,
    new_G3007gat, new_G3010gat, new_G3014gat, new_G3015gat, new_G3016gat,
    new_G3019gat, new_G3022gat, new_G3026gat, new_G3027gat, new_G3028gat,
    new_G3031gat, new_G3034gat, new_G3037gat, new_G3040gat, new_G3043gat,
    new_G3046gat, new_G3049gat, new_G3052gat, new_G3055gat, new_G3058gat,
    new_G3062gat, new_G3063gat, new_G3064gat, new_G3067gat, new_G3070gat,
    new_G3074gat, new_G3075gat, new_G3076gat, new_G3079gat, new_G3083gat,
    new_G3087gat, new_G3091gat, new_G3095gat, new_G3099gat, new_G3103gat,
    new_G3107gat, new_G3111gat, new_G3115gat, new_G3119gat, new_G3120gat,
    new_G3121gat, new_G3124gat, new_G3127gat, new_G3131gat, new_G3132gat,
    new_G3133gat, new_G3136gat, new_G3140gat, new_G3141gat, new_G3142gat,
    new_G3145gat, new_G3146gat, new_G3147gat, new_G3150gat, new_G3151gat,
    new_G3152gat, new_G3155gat, new_G3156gat, new_G3157gat, new_G3160gat,
    new_G3161gat, new_G3162gat, new_G3165gat, new_G3166gat, new_G3167gat,
    new_G3170gat, new_G3171gat, new_G3172gat, new_G3175gat, new_G3176gat,
    new_G3177gat, new_G3180gat, new_G3181gat, new_G3182gat, new_G3185gat,
    new_G3186gat, new_G3187gat, new_G3190gat, new_G3193gat, new_G3197gat,
    new_G3198gat, new_G3199gat, new_G3202gat, new_G3206gat, new_G3207gat,
    new_G3208gat, new_G3212gat, new_G3215gat, new_G3218gat, new_G3221gat,
    new_G3224gat, new_G3227gat, new_G3230gat, new_G3233gat, new_G3236gat,
    new_G3239gat, new_G3243gat, new_G3244gat, new_G3245gat, new_G3248gat,
    new_G3252gat, new_G3253gat, new_G3254gat, new_G3257gat, new_G3260gat,
    new_G3264gat, new_G3268gat, new_G3272gat, new_G3276gat, new_G3280gat,
    new_G3284gat, new_G3288gat, new_G3292gat, new_G3296gat, new_G3300gat,
    new_G3301gat, new_G3302gat, new_G3305gat, new_G3309gat, new_G3310gat,
    new_G3311gat, new_G3314gat, new_G3317gat, new_G3321gat, new_G3322gat,
    new_G3323gat, new_G3324gat, new_G3325gat, new_G3326gat, new_G3327gat,
    new_G3328gat, new_G3329gat, new_G3330gat, new_G3331gat, new_G3332gat,
    new_G3333gat, new_G3334gat, new_G3335gat, new_G3336gat, new_G3337gat,
    new_G3338gat, new_G3339gat, new_G3340gat, new_G3341gat, new_G3344gat,
    new_G3348gat, new_G3349gat, new_G3350gat, new_G3353gat, new_G3356gat,
    new_G3360gat, new_G3361gat, new_G3362gat, new_G3365gat, new_G3368gat,
    new_G3371gat, new_G3374gat, new_G3377gat, new_G3380gat, new_G3383gat,
    new_G3386gat, new_G3389gat, new_G3392gat, new_G3396gat, new_G3397gat,
    new_G3398gat, new_G3401gat, new_G3404gat, new_G3408gat, new_G3409gat,
    new_G3410gat, new_G3413gat, new_G3417gat, new_G3421gat, new_G3425gat,
    new_G3429gat, new_G3433gat, new_G3437gat, new_G3441gat, new_G3445gat,
    new_G3449gat, new_G3453gat, new_G3454gat, new_G3455gat, new_G3458gat,
    new_G3461gat, new_G3465gat, new_G3466gat, new_G3467gat, new_G3470gat,
    new_G3474gat, new_G3475gat, new_G3476gat, new_G3479gat, new_G3480gat,
    new_G3481gat, new_G3484gat, new_G3485gat, new_G3486gat, new_G3489gat,
    new_G3490gat, new_G3491gat, new_G3494gat, new_G3495gat, new_G3496gat,
    new_G3499gat, new_G3500gat, new_G3501gat, new_G3504gat, new_G3505gat,
    new_G3506gat, new_G3509gat, new_G3510gat, new_G3511gat, new_G3514gat,
    new_G3515gat, new_G3516gat, new_G3519gat, new_G3520gat, new_G3521gat,
    new_G3524gat, new_G3527gat, new_G3531gat, new_G3532gat, new_G3533gat,
    new_G3536gat, new_G3540gat, new_G3541gat, new_G3542gat, new_G3545gat,
    new_G3548gat, new_G3553gat, new_G3556gat, new_G3559gat, new_G3562gat,
    new_G3565gat, new_G3568gat, new_G3571gat, new_G3574gat, new_G3577gat,
    new_G3581gat, new_G3582gat, new_G3583gat, new_G3586gat, new_G3590gat,
    new_G3591gat, new_G3592gat, new_G3595gat, new_G3598gat, new_G3602gat,
    new_G3603gat, new_G3604gat, new_G3608gat, new_G3612gat, new_G3616gat,
    new_G3620gat, new_G3624gat, new_G3628gat, new_G3632gat, new_G3636gat,
    new_G3637gat, new_G3638gat, new_G3641gat, new_G3645gat, new_G3646gat,
    new_G3647gat, new_G3650gat, new_G3653gat, new_G3657gat, new_G3658gat,
    new_G3659gat, new_G3662gat, new_G3663gat, new_G3664gat, new_G3665gat,
    new_G3666gat, new_G3667gat, new_G3668gat, new_G3669gat, new_G3670gat,
    new_G3671gat, new_G3672gat, new_G3673gat, new_G3674gat, new_G3675gat,
    new_G3676gat, new_G3677gat, new_G3678gat, new_G3681gat, new_G3685gat,
    new_G3686gat, new_G3687gat, new_G3690gat, new_G3693gat, new_G3697gat,
    new_G3698gat, new_G3699gat, new_G3702gat, new_G3706gat, new_G3709gat,
    new_G3712gat, new_G3715gat, new_G3718gat, new_G3721gat, new_G3724gat,
    new_G3727gat, new_G3730gat, new_G3734gat, new_G3735gat, new_G3736gat,
    new_G3739gat, new_G3742gat, new_G3746gat, new_G3747gat, new_G3748gat,
    new_G3751gat, new_G3755gat, new_G3756gat, new_G3757gat, new_G3760gat,
    new_G3764gat, new_G3768gat, new_G3772gat, new_G3776gat, new_G3780gat,
    new_G3784gat, new_G3788gat, new_G3792gat, new_G3793gat, new_G3794gat,
    new_G3797gat, new_G3800gat, new_G3804gat, new_G3805gat, new_G3806gat,
    new_G3809gat, new_G3813gat, new_G3814gat, new_G3815gat, new_G3818gat,
    new_G3821gat, new_G3825gat, new_G3826gat, new_G3827gat, new_G3830gat,
    new_G3831gat, new_G3832gat, new_G3835gat, new_G3836gat, new_G3837gat,
    new_G3840gat, new_G3841gat, new_G3842gat, new_G3845gat, new_G3846gat,
    new_G3847gat, new_G3850gat, new_G3851gat, new_G3852gat, new_G3855gat,
    new_G3856gat, new_G3857gat, new_G3860gat, new_G3861gat, new_G3862gat,
    new_G3865gat, new_G3868gat, new_G3872gat, new_G3873gat, new_G3874gat,
    new_G3877gat, new_G3881gat, new_G3882gat, new_G3883gat, new_G3886gat,
    new_G3889gat, new_G3893gat, new_G3894gat, new_G3896gat, new_G3899gat,
    new_G3902gat, new_G3905gat, new_G3908gat, new_G3911gat, new_G3914gat,
    new_G3917gat, new_G3921gat, new_G3922gat, new_G3923gat, new_G3926gat,
    new_G3930gat, new_G3931gat, new_G3932gat, new_G3935gat, new_G3938gat,
    new_G3942gat, new_G3943gat, new_G3944gat, new_G3947gat, new_G3951gat,
    new_G3955gat, new_G3959gat, new_G3963gat, new_G3967gat, new_G3971gat,
    new_G3975gat, new_G3976gat, new_G3977gat, new_G3980gat, new_G3984gat,
    new_G3985gat, new_G3986gat, new_G3989gat, new_G3992gat, new_G3996gat,
    new_G3997gat, new_G3998gat, new_G4001gat, new_G4005gat, new_G4006gat,
    new_G4007gat, new_G4008gat, new_G4009gat, new_G4010gat, new_G4011gat,
    new_G4012gat, new_G4013gat, new_G4014gat, new_G4015gat, new_G4016gat,
    new_G4017gat, new_G4018gat, new_G4019gat, new_G4022gat, new_G4026gat,
    new_G4027gat, new_G4028gat, new_G4031gat, new_G4034gat, new_G4038gat,
    new_G4039gat, new_G4040gat, new_G4043gat, new_G4047gat, new_G4048gat,
    new_G4049gat, new_G4052gat, new_G4055gat, new_G4058gat, new_G4061gat,
    new_G4064gat, new_G4067gat, new_G4070gat, new_G4073gat, new_G4077gat,
    new_G4078gat, new_G4079gat, new_G4082gat, new_G4085gat, new_G4089gat,
    new_G4090gat, new_G4091gat, new_G4094gat, new_G4098gat, new_G4099gat,
    new_G4100gat, new_G4103gat, new_G4106gat, new_G4110gat, new_G4114gat,
    new_G4118gat, new_G4122gat, new_G4126gat, new_G4130gat, new_G4134gat,
    new_G4138gat, new_G4139gat, new_G4140gat, new_G4143gat, new_G4146gat,
    new_G4150gat, new_G4151gat, new_G4152gat, new_G4155gat, new_G4159gat,
    new_G4160gat, new_G4161gat, new_G4164gat, new_G4167gat, new_G4171gat,
    new_G4172gat, new_G4173gat, new_G4174gat, new_G4175gat, new_G4178gat,
    new_G4179gat, new_G4180gat, new_G4183gat, new_G4184gat, new_G4185gat,
    new_G4188gat, new_G4189gat, new_G4190gat, new_G4193gat, new_G4194gat,
    new_G4195gat, new_G4198gat, new_G4199gat, new_G4200gat, new_G4203gat,
    new_G4204gat, new_G4205gat, new_G4208gat, new_G4211gat, new_G4215gat,
    new_G4216gat, new_G4217gat, new_G4220gat, new_G4224gat, new_G4225gat,
    new_G4226gat, new_G4229gat, new_G4232gat, new_G4236gat, new_G4237gat,
    new_G4238gat, new_G4242gat, new_G4245gat, new_G4248gat, new_G4251gat,
    new_G4254gat, new_G4257gat, new_G4260gat, new_G4264gat, new_G4265gat,
    new_G4266gat, new_G4269gat, new_G4273gat, new_G4274gat, new_G4275gat,
    new_G4278gat, new_G4281gat, new_G4285gat, new_G4286gat, new_G4287gat,
    new_G4290gat, new_G4294gat, new_G4298gat, new_G4302gat, new_G4306gat,
    new_G4310gat, new_G4314gat, new_G4318gat, new_G4319gat, new_G4320gat,
    new_G4323gat, new_G4327gat, new_G4328gat, new_G4329gat, new_G4332gat,
    new_G4335gat, new_G4339gat, new_G4340gat, new_G4341gat, new_G4344gat,
    new_G4348gat, new_G4349gat, new_G4350gat, new_G4353gat, new_G4354gat,
    new_G4355gat, new_G4356gat, new_G4357gat, new_G4358gat, new_G4359gat,
    new_G4360gat, new_G4361gat, new_G4362gat, new_G4363gat, new_G4364gat,
    new_G4365gat, new_G4368gat, new_G4372gat, new_G4373gat, new_G4374gat,
    new_G4377gat, new_G4380gat, new_G4384gat, new_G4385gat, new_G4386gat,
    new_G4389gat, new_G4393gat, new_G4394gat, new_G4395gat, new_G4398gat,
    new_G4401gat, new_G4405gat, new_G4408gat, new_G4411gat, new_G4414gat,
    new_G4417gat, new_G4420gat, new_G4423gat, new_G4427gat, new_G4428gat,
    new_G4429gat, new_G4432gat, new_G4435gat, new_G4439gat, new_G4440gat,
    new_G4441gat, new_G4444gat, new_G4448gat, new_G4449gat, new_G4450gat,
    new_G4453gat, new_G4456gat, new_G4460gat, new_G4461gat, new_G4462gat,
    new_G4466gat, new_G4470gat, new_G4474gat, new_G4478gat, new_G4482gat,
    new_G4486gat, new_G4487gat, new_G4488gat, new_G4491gat, new_G4494gat,
    new_G4498gat, new_G4499gat, new_G4500gat, new_G4503gat, new_G4507gat,
    new_G4508gat, new_G4509gat, new_G4512gat, new_G4515gat, new_G4519gat,
    new_G4520gat, new_G4521gat, new_G4524gat, new_G4525gat, new_G4526gat,
    new_G4529gat, new_G4530gat, new_G4531gat, new_G4534gat, new_G4535gat,
    new_G4536gat, new_G4539gat, new_G4540gat, new_G4541gat, new_G4544gat,
    new_G4545gat, new_G4546gat, new_G4549gat, new_G4550gat, new_G4551gat,
    new_G4554gat, new_G4557gat, new_G4561gat, new_G4562gat, new_G4563gat,
    new_G4566gat, new_G4570gat, new_G4571gat, new_G4572gat, new_G4575gat,
    new_G4578gat, new_G4582gat, new_G4583gat, new_G4584gat, new_G4587gat,
    new_G4592gat, new_G4595gat, new_G4598gat, new_G4601gat, new_G4604gat,
    new_G4607gat, new_G4611gat, new_G4612gat, new_G4613gat, new_G4616gat,
    new_G4620gat, new_G4621gat, new_G4622gat, new_G4625gat, new_G4628gat,
    new_G4632gat, new_G4633gat, new_G4634gat, new_G4637gat, new_G4641gat,
    new_G4642gat, new_G4643gat, new_G4646gat, new_G4650gat, new_G4654gat,
    new_G4658gat, new_G4662gat, new_G4666gat, new_G4667gat, new_G4668gat,
    new_G4671gat, new_G4675gat, new_G4676gat, new_G4677gat, new_G4680gat,
    new_G4683gat, new_G4687gat, new_G4688gat, new_G4689gat, new_G4692gat,
    new_G4696gat, new_G4697gat, new_G4698gat, new_G4701gat, new_G4704gat,
    new_G4708gat, new_G4709gat, new_G4710gat, new_G4711gat, new_G4712gat,
    new_G4713gat, new_G4714gat, new_G4715gat, new_G4716gat, new_G4717gat,
    new_G4718gat, new_G4721gat, new_G4725gat, new_G4726gat, new_G4727gat,
    new_G4730gat, new_G4733gat, new_G4737gat, new_G4738gat, new_G4739gat,
    new_G4742gat, new_G4746gat, new_G4747gat, new_G4748gat, new_G4751gat,
    new_G4754gat, new_G4758gat, new_G4759gat, new_G4760gat, new_G4763gat,
    new_G4766gat, new_G4769gat, new_G4772gat, new_G4775gat, new_G4779gat,
    new_G4780gat, new_G4781gat, new_G4784gat, new_G4787gat, new_G4791gat,
    new_G4792gat, new_G4793gat, new_G4796gat, new_G4800gat, new_G4801gat,
    new_G4802gat, new_G4805gat, new_G4808gat, new_G4812gat, new_G4813gat,
    new_G4814gat, new_G4817gat, new_G4821gat, new_G4825gat, new_G4829gat,
    new_G4833gat, new_G4837gat, new_G4838gat, new_G4839gat, new_G4842gat,
    new_G4845gat, new_G4849gat, new_G4850gat, new_G4851gat, new_G4854gat,
    new_G4858gat, new_G4859gat, new_G4860gat, new_G4863gat, new_G4866gat,
    new_G4870gat, new_G4871gat, new_G4872gat, new_G4875gat, new_G4879gat,
    new_G4880gat, new_G4881gat, new_G4884gat, new_G4885gat, new_G4886gat,
    new_G4889gat, new_G4890gat, new_G4891gat, new_G4894gat, new_G4895gat,
    new_G4896gat, new_G4899gat, new_G4900gat, new_G4901gat, new_G4904gat,
    new_G4907gat, new_G4911gat, new_G4912gat, new_G4913gat, new_G4916gat,
    new_G4920gat, new_G4921gat, new_G4922gat, new_G4925gat, new_G4928gat,
    new_G4932gat, new_G4933gat, new_G4934gat, new_G4937gat, new_G4941gat,
    new_G4942gat, new_G4943gat, new_G4947gat, new_G4950gat, new_G4953gat,
    new_G4956gat, new_G4959gat, new_G4963gat, new_G4964gat, new_G4965gat,
    new_G4968gat, new_G4972gat, new_G4973gat, new_G4974gat, new_G4977gat,
    new_G4980gat, new_G4984gat, new_G4985gat, new_G4986gat, new_G4989gat,
    new_G4993gat, new_G4994gat, new_G4995gat, new_G4998gat, new_G5001gat,
    new_G5005gat, new_G5009gat, new_G5013gat, new_G5017gat, new_G5021gat,
    new_G5022gat, new_G5023gat, new_G5026gat, new_G5030gat, new_G5031gat,
    new_G5032gat, new_G5035gat, new_G5038gat, new_G5042gat, new_G5043gat,
    new_G5044gat, new_G5047gat, new_G5051gat, new_G5052gat, new_G5053gat,
    new_G5056gat, new_G5059gat, new_G5063gat, new_G5064gat, new_G5065gat,
    new_G5066gat, new_G5067gat, new_G5068gat, new_G5069gat, new_G5070gat,
    new_G5071gat, new_G5072gat, new_G5073gat, new_G5076gat, new_G5080gat,
    new_G5081gat, new_G5082gat, new_G5085gat, new_G5088gat, new_G5092gat,
    new_G5093gat, new_G5094gat, new_G5097gat, new_G5101gat, new_G5102gat,
    new_G5103gat, new_G5106gat, new_G5109gat, new_G5113gat, new_G5114gat,
    new_G5115gat, new_G5118gat, new_G5121gat, new_G5124gat, new_G5127gat,
    new_G5130gat, new_G5134gat, new_G5135gat, new_G5136gat, new_G5139gat,
    new_G5142gat, new_G5146gat, new_G5147gat, new_G5148gat, new_G5151gat,
    new_G5155gat, new_G5156gat, new_G5157gat, new_G5160gat, new_G5163gat,
    new_G5167gat, new_G5168gat, new_G5169gat, new_G5172gat, new_G5176gat,
    new_G5180gat, new_G5184gat, new_G5188gat, new_G5192gat, new_G5193gat,
    new_G5194gat, new_G5197gat, new_G5200gat, new_G5204gat, new_G5205gat,
    new_G5206gat, new_G5209gat, new_G5213gat, new_G5214gat, new_G5215gat,
    new_G5218gat, new_G5221gat, new_G5225gat, new_G5226gat, new_G5227gat,
    new_G5230gat, new_G5234gat, new_G5235gat, new_G5236gat, new_G5239gat,
    new_G5240gat, new_G5241gat, new_G5244gat, new_G5245gat, new_G5246gat,
    new_G5249gat, new_G5250gat, new_G5251gat, new_G5254gat, new_G5255gat,
    new_G5256gat, new_G5259gat, new_G5262gat, new_G5266gat, new_G5267gat,
    new_G5268gat, new_G5271gat, new_G5275gat, new_G5276gat, new_G5277gat,
    new_G5280gat, new_G5283gat, new_G5287gat, new_G5288gat, new_G5289gat,
    new_G5292gat, new_G5296gat, new_G5297gat, new_G5298gat, new_G5301gat,
    new_G5304gat, new_G5309gat, new_G5312gat, new_G5315gat, new_G5318gat,
    new_G5322gat, new_G5323gat, new_G5324gat, new_G5327gat, new_G5331gat,
    new_G5332gat, new_G5333gat, new_G5336gat, new_G5339gat, new_G5343gat,
    new_G5344gat, new_G5345gat, new_G5348gat, new_G5352gat, new_G5353gat,
    new_G5354gat, new_G5357gat, new_G5360gat, new_G5364gat, new_G5365gat,
    new_G5366gat, new_G5370gat, new_G5374gat, new_G5378gat, new_G5379gat,
    new_G5380gat, new_G5383gat, new_G5387gat, new_G5388gat, new_G5389gat,
    new_G5392gat, new_G5395gat, new_G5399gat, new_G5400gat, new_G5401gat,
    new_G5404gat, new_G5408gat, new_G5409gat, new_G5410gat, new_G5413gat,
    new_G5416gat, new_G5420gat, new_G5421gat, new_G5422gat, new_G5425gat,
    new_G5426gat, new_G5427gat, new_G5428gat, new_G5429gat, new_G5430gat,
    new_G5431gat, new_G5434gat, new_G5438gat, new_G5439gat, new_G5440gat,
    new_G5443gat, new_G5446gat, new_G5450gat, new_G5451gat, new_G5452gat,
    new_G5455gat, new_G5459gat, new_G5460gat, new_G5461gat, new_G5464gat,
    new_G5467gat, new_G5471gat, new_G5472gat, new_G5473gat, new_G5476gat,
    new_G5480gat, new_G5483gat, new_G5486gat, new_G5489gat, new_G5493gat,
    new_G5494gat, new_G5495gat, new_G5498gat, new_G5501gat, new_G5505gat,
    new_G5506gat, new_G5507gat, new_G5510gat, new_G5514gat, new_G5515gat,
    new_G5516gat, new_G5519gat, new_G5522gat, new_G5526gat, new_G5527gat,
    new_G5528gat, new_G5531gat, new_G5535gat, new_G5536gat, new_G5537gat,
    new_G5540gat, new_G5544gat, new_G5548gat, new_G5552gat, new_G5553gat,
    new_G5554gat, new_G5557gat, new_G5560gat, new_G5564gat, new_G5565gat,
    new_G5566gat, new_G5569gat, new_G5573gat, new_G5574gat, new_G5575gat,
    new_G5578gat, new_G5581gat, new_G5585gat, new_G5586gat, new_G5587gat,
    new_G5590gat, new_G5594gat, new_G5595gat, new_G5596gat, new_G5599gat,
    new_G5602gat, new_G5606gat, new_G5607gat, new_G5608gat, new_G5611gat,
    new_G5612gat, new_G5613gat, new_G5616gat, new_G5617gat, new_G5618gat,
    new_G5621gat, new_G5624gat, new_G5628gat, new_G5629gat, new_G5630gat,
    new_G5633gat, new_G5637gat, new_G5638gat, new_G5639gat, new_G5642gat,
    new_G5645gat, new_G5649gat, new_G5650gat, new_G5651gat, new_G5654gat,
    new_G5658gat, new_G5659gat, new_G5660gat, new_G5663gat, new_G5666gat,
    new_G5670gat, new_G5671gat, new_G5673gat, new_G5676gat, new_G5679gat,
    new_G5683gat, new_G5684gat, new_G5685gat, new_G5688gat, new_G5692gat,
    new_G5693gat, new_G5694gat, new_G5697gat, new_G5700gat, new_G5704gat,
    new_G5705gat, new_G5706gat, new_G5709gat, new_G5713gat, new_G5714gat,
    new_G5715gat, new_G5718gat, new_G5721gat, new_G5725gat, new_G5726gat,
    new_G5727gat, new_G5730gat, new_G5734gat, new_G5738gat, new_G5739gat,
    new_G5740gat, new_G5743gat, new_G5747gat, new_G5748gat, new_G5749gat,
    new_G5752gat, new_G5755gat, new_G5759gat, new_G5760gat, new_G5761gat,
    new_G5764gat, new_G5768gat, new_G5769gat, new_G5770gat, new_G5773gat,
    new_G5776gat, new_G5780gat, new_G5781gat, new_G5782gat, new_G5785gat,
    new_G5786gat, new_G5787gat, new_G5788gat, new_G5789gat, new_G5792gat,
    new_G5796gat, new_G5797gat, new_G5798gat, new_G5801gat, new_G5804gat,
    new_G5808gat, new_G5809gat, new_G5810gat, new_G5813gat, new_G5817gat,
    new_G5818gat, new_G5819gat, new_G5822gat, new_G5825gat, new_G5829gat,
    new_G5830gat, new_G5831gat, new_G5834gat, new_G5837gat, new_G5840gat,
    new_G5844gat, new_G5845gat, new_G5846gat, new_G5849gat, new_G5852gat,
    new_G5856gat, new_G5857gat, new_G5858gat, new_G5861gat, new_G5865gat,
    new_G5866gat, new_G5867gat, new_G5870gat, new_G5873gat, new_G5877gat,
    new_G5878gat, new_G5879gat, new_G5882gat, new_G5886gat, new_G5890gat,
    new_G5891gat, new_G5892gat, new_G5895gat, new_G5898gat, new_G5902gat,
    new_G5903gat, new_G5904gat, new_G5907gat, new_G5911gat, new_G5912gat,
    new_G5913gat, new_G5916gat, new_G5919gat, new_G5923gat, new_G5924gat,
    new_G5925gat, new_G5928gat, new_G5929gat, new_G5930gat, new_G5933gat,
    new_G5934gat, new_G5935gat, new_G5938gat, new_G5941gat, new_G5945gat,
    new_G5946gat, new_G5947gat, new_G5950gat, new_G5954gat, new_G5955gat,
    new_G5956gat, new_G5959gat, new_G5962gat, new_G5966gat, new_G5967gat,
    new_G5968gat, new_G5972gat, new_G5975gat, new_G5979gat, new_G5980gat,
    new_G5981gat, new_G5984gat, new_G5988gat, new_G5989gat, new_G5990gat,
    new_G5993gat, new_G5996gat, new_G6000gat, new_G6001gat, new_G6002gat,
    new_G6005gat, new_G6009gat, new_G6010gat, new_G6011gat, new_G6014gat,
    new_G6018gat, new_G6019gat, new_G6020gat, new_G6023gat, new_G6026gat,
    new_G6030gat, new_G6031gat, new_G6032gat, new_G6035gat, new_G6036gat,
    new_G6037gat, new_G6040gat, new_G6044gat, new_G6045gat, new_G6046gat,
    new_G6049gat, new_G6052gat, new_G6056gat, new_G6057gat, new_G6058gat,
    new_G6061gat, new_G6064gat, new_G6068gat, new_G6069gat, new_G6070gat,
    new_G6073gat, new_G6076gat, new_G6080gat, new_G6081gat, new_G6082gat,
    new_G6085gat, new_G6089gat, new_G6090gat, new_G6091gat, new_G6094gat,
    new_G6097gat, new_G6101gat, new_G6102gat, new_G6103gat, new_G6106gat,
    new_G6107gat, new_G6108gat, new_G6111gat, new_G6114gat, new_G6118gat,
    new_G6119gat, new_G6120gat, new_G6124gat, new_G6128gat, new_G6129gat,
    new_G6130gat, new_G6133gat, new_G6134gat, new_G6135gat, new_G6138gat,
    new_G6141gat, new_G6145gat, new_G6146gat, new_G6147gat, new_G6151gat,
    new_G6155gat, new_G6156gat, new_G6157gat, new_G6161gat, new_G6165gat,
    new_G6166gat, new_G6167gat, new_G6171gat, new_G6175gat, new_G6176gat,
    new_G6177gat, new_G6181gat, new_G6185gat, new_G6186gat, new_G6187gat,
    new_G6191gat, new_G6195gat, new_G6196gat, new_G6197gat, new_G6201gat,
    new_G6205gat, new_G6206gat, new_G6207gat, new_G6211gat, new_G6215gat,
    new_G6216gat, new_G6217gat, new_G6221gat, new_G6225gat, new_G6226gat,
    new_G6227gat, new_G6231gat, new_G6235gat, new_G6236gat, new_G6237gat,
    new_G6241gat, new_G6245gat, new_G6246gat, new_G6247gat, new_G6251gat,
    new_G6255gat, new_G6256gat, new_G6257gat, new_G6261gat, new_G6265gat,
    new_G6266gat, new_G6267gat, new_G6271gat, new_G6275gat, new_G6276gat,
    new_G6277gat, new_G6281gat, new_G6285gat, new_G6286gat;
  assign G545gat = G1gat & G273gat;
  assign new_G546gat = G1gat & G290gat;
  assign new_G549gat = G1gat & G307gat;
  assign new_G552gat = G1gat & G324gat;
  assign new_G555gat = G1gat & G341gat;
  assign new_G558gat = G1gat & G358gat;
  assign new_G561gat = G1gat & G375gat;
  assign new_G564gat = G1gat & G392gat;
  assign new_G567gat = G1gat & G409gat;
  assign new_G570gat = G1gat & G426gat;
  assign new_G573gat = G1gat & G443gat;
  assign new_G576gat = G1gat & G460gat;
  assign new_G579gat = G1gat & G477gat;
  assign new_G582gat = G1gat & G494gat;
  assign new_G585gat = G1gat & G511gat;
  assign new_G588gat = G1gat & G528gat;
  assign new_G591gat = G18gat & G273gat;
  assign new_G594gat = G18gat & G290gat;
  assign new_G597gat = G18gat & G307gat;
  assign new_G600gat = G18gat & G324gat;
  assign new_G603gat = G18gat & G341gat;
  assign new_G606gat = G18gat & G358gat;
  assign new_G609gat = G18gat & G375gat;
  assign new_G612gat = G18gat & G392gat;
  assign new_G615gat = G18gat & G409gat;
  assign new_G618gat = G18gat & G426gat;
  assign new_G621gat = G18gat & G443gat;
  assign new_G624gat = G18gat & G460gat;
  assign new_G627gat = G18gat & G477gat;
  assign new_G630gat = G18gat & G494gat;
  assign new_G633gat = G18gat & G511gat;
  assign new_G636gat = G18gat & G528gat;
  assign new_G639gat = G35gat & G273gat;
  assign new_G642gat = G35gat & G290gat;
  assign new_G645gat = G35gat & G307gat;
  assign new_G648gat = G35gat & G324gat;
  assign new_G651gat = G35gat & G341gat;
  assign new_G654gat = G35gat & G358gat;
  assign new_G657gat = G35gat & G375gat;
  assign new_G660gat = G35gat & G392gat;
  assign new_G663gat = G35gat & G409gat;
  assign new_G666gat = G35gat & G426gat;
  assign new_G669gat = G35gat & G443gat;
  assign new_G672gat = G35gat & G460gat;
  assign new_G675gat = G35gat & G477gat;
  assign new_G678gat = G35gat & G494gat;
  assign new_G681gat = G35gat & G511gat;
  assign new_G684gat = G35gat & G528gat;
  assign new_G687gat = G52gat & G273gat;
  assign new_G690gat = G52gat & G290gat;
  assign new_G693gat = G52gat & G307gat;
  assign new_G696gat = G52gat & G324gat;
  assign new_G699gat = G52gat & G341gat;
  assign new_G702gat = G52gat & G358gat;
  assign new_G705gat = G52gat & G375gat;
  assign new_G708gat = G52gat & G392gat;
  assign new_G711gat = G52gat & G409gat;
  assign new_G714gat = G52gat & G426gat;
  assign new_G717gat = G52gat & G443gat;
  assign new_G720gat = G52gat & G460gat;
  assign new_G723gat = G52gat & G477gat;
  assign new_G726gat = G52gat & G494gat;
  assign new_G729gat = G52gat & G511gat;
  assign new_G732gat = G52gat & G528gat;
  assign new_G735gat = G69gat & G273gat;
  assign new_G738gat = G69gat & G290gat;
  assign new_G741gat = G69gat & G307gat;
  assign new_G744gat = G69gat & G324gat;
  assign new_G747gat = G69gat & G341gat;
  assign new_G750gat = G69gat & G358gat;
  assign new_G753gat = G69gat & G375gat;
  assign new_G756gat = G69gat & G392gat;
  assign new_G759gat = G69gat & G409gat;
  assign new_G762gat = G69gat & G426gat;
  assign new_G765gat = G69gat & G443gat;
  assign new_G768gat = G69gat & G460gat;
  assign new_G771gat = G69gat & G477gat;
  assign new_G774gat = G69gat & G494gat;
  assign new_G777gat = G69gat & G511gat;
  assign new_G780gat = G69gat & G528gat;
  assign new_G783gat = G86gat & G273gat;
  assign new_G786gat = G86gat & G290gat;
  assign new_G789gat = G86gat & G307gat;
  assign new_G792gat = G86gat & G324gat;
  assign new_G795gat = G86gat & G341gat;
  assign new_G798gat = G86gat & G358gat;
  assign new_G801gat = G86gat & G375gat;
  assign new_G804gat = G86gat & G392gat;
  assign new_G807gat = G86gat & G409gat;
  assign new_G810gat = G86gat & G426gat;
  assign new_G813gat = G86gat & G443gat;
  assign new_G816gat = G86gat & G460gat;
  assign new_G819gat = G86gat & G477gat;
  assign new_G822gat = G86gat & G494gat;
  assign new_G825gat = G86gat & G511gat;
  assign new_G828gat = G86gat & G528gat;
  assign new_G831gat = G103gat & G273gat;
  assign new_G834gat = G103gat & G290gat;
  assign new_G837gat = G103gat & G307gat;
  assign new_G840gat = G103gat & G324gat;
  assign new_G843gat = G103gat & G341gat;
  assign new_G846gat = G103gat & G358gat;
  assign new_G849gat = G103gat & G375gat;
  assign new_G852gat = G103gat & G392gat;
  assign new_G855gat = G103gat & G409gat;
  assign new_G858gat = G103gat & G426gat;
  assign new_G861gat = G103gat & G443gat;
  assign new_G864gat = G103gat & G460gat;
  assign new_G867gat = G103gat & G477gat;
  assign new_G870gat = G103gat & G494gat;
  assign new_G873gat = G103gat & G511gat;
  assign new_G876gat = G103gat & G528gat;
  assign new_G879gat = G120gat & G273gat;
  assign new_G882gat = G120gat & G290gat;
  assign new_G885gat = G120gat & G307gat;
  assign new_G888gat = G120gat & G324gat;
  assign new_G891gat = G120gat & G341gat;
  assign new_G894gat = G120gat & G358gat;
  assign new_G897gat = G120gat & G375gat;
  assign new_G900gat = G120gat & G392gat;
  assign new_G903gat = G120gat & G409gat;
  assign new_G906gat = G120gat & G426gat;
  assign new_G909gat = G120gat & G443gat;
  assign new_G912gat = G120gat & G460gat;
  assign new_G915gat = G120gat & G477gat;
  assign new_G918gat = G120gat & G494gat;
  assign new_G921gat = G120gat & G511gat;
  assign new_G924gat = G120gat & G528gat;
  assign new_G927gat = G137gat & G273gat;
  assign new_G930gat = G137gat & G290gat;
  assign new_G933gat = G137gat & G307gat;
  assign new_G936gat = G137gat & G324gat;
  assign new_G939gat = G137gat & G341gat;
  assign new_G942gat = G137gat & G358gat;
  assign new_G945gat = G137gat & G375gat;
  assign new_G948gat = G137gat & G392gat;
  assign new_G951gat = G137gat & G409gat;
  assign new_G954gat = G137gat & G426gat;
  assign new_G957gat = G137gat & G443gat;
  assign new_G960gat = G137gat & G460gat;
  assign new_G963gat = G137gat & G477gat;
  assign new_G966gat = G137gat & G494gat;
  assign new_G969gat = G137gat & G511gat;
  assign new_G972gat = G137gat & G528gat;
  assign new_G975gat = G154gat & G273gat;
  assign new_G978gat = G154gat & G290gat;
  assign new_G981gat = G154gat & G307gat;
  assign new_G984gat = G154gat & G324gat;
  assign new_G987gat = G154gat & G341gat;
  assign new_G990gat = G154gat & G358gat;
  assign new_G993gat = G154gat & G375gat;
  assign new_G996gat = G154gat & G392gat;
  assign new_G999gat = G154gat & G409gat;
  assign new_G1002gat = G154gat & G426gat;
  assign new_G1005gat = G154gat & G443gat;
  assign new_G1008gat = G154gat & G460gat;
  assign new_G1011gat = G154gat & G477gat;
  assign new_G1014gat = G154gat & G494gat;
  assign new_G1017gat = G154gat & G511gat;
  assign new_G1020gat = G154gat & G528gat;
  assign new_G1023gat = G171gat & G273gat;
  assign new_G1026gat = G171gat & G290gat;
  assign new_G1029gat = G171gat & G307gat;
  assign new_G1032gat = G171gat & G324gat;
  assign new_G1035gat = G171gat & G341gat;
  assign new_G1038gat = G171gat & G358gat;
  assign new_G1041gat = G171gat & G375gat;
  assign new_G1044gat = G171gat & G392gat;
  assign new_G1047gat = G171gat & G409gat;
  assign new_G1050gat = G171gat & G426gat;
  assign new_G1053gat = G171gat & G443gat;
  assign new_G1056gat = G171gat & G460gat;
  assign new_G1059gat = G171gat & G477gat;
  assign new_G1062gat = G171gat & G494gat;
  assign new_G1065gat = G171gat & G511gat;
  assign new_G1068gat = G171gat & G528gat;
  assign new_G1071gat = G188gat & G273gat;
  assign new_G1074gat = G188gat & G290gat;
  assign new_G1077gat = G188gat & G307gat;
  assign new_G1080gat = G188gat & G324gat;
  assign new_G1083gat = G188gat & G341gat;
  assign new_G1086gat = G188gat & G358gat;
  assign new_G1089gat = G188gat & G375gat;
  assign new_G1092gat = G188gat & G392gat;
  assign new_G1095gat = G188gat & G409gat;
  assign new_G1098gat = G188gat & G426gat;
  assign new_G1101gat = G188gat & G443gat;
  assign new_G1104gat = G188gat & G460gat;
  assign new_G1107gat = G188gat & G477gat;
  assign new_G1110gat = G188gat & G494gat;
  assign new_G1113gat = G188gat & G511gat;
  assign new_G1116gat = G188gat & G528gat;
  assign new_G1119gat = G205gat & G273gat;
  assign new_G1122gat = G205gat & G290gat;
  assign new_G1125gat = G205gat & G307gat;
  assign new_G1128gat = G205gat & G324gat;
  assign new_G1131gat = G205gat & G341gat;
  assign new_G1134gat = G205gat & G358gat;
  assign new_G1137gat = G205gat & G375gat;
  assign new_G1140gat = G205gat & G392gat;
  assign new_G1143gat = G205gat & G409gat;
  assign new_G1146gat = G205gat & G426gat;
  assign new_G1149gat = G205gat & G443gat;
  assign new_G1152gat = G205gat & G460gat;
  assign new_G1155gat = G205gat & G477gat;
  assign new_G1158gat = G205gat & G494gat;
  assign new_G1161gat = G205gat & G511gat;
  assign new_G1164gat = G205gat & G528gat;
  assign new_G1167gat = G222gat & G273gat;
  assign new_G1170gat = G222gat & G290gat;
  assign new_G1173gat = G222gat & G307gat;
  assign new_G1176gat = G222gat & G324gat;
  assign new_G1179gat = G222gat & G341gat;
  assign new_G1182gat = G222gat & G358gat;
  assign new_G1185gat = G222gat & G375gat;
  assign new_G1188gat = G222gat & G392gat;
  assign new_G1191gat = G222gat & G409gat;
  assign new_G1194gat = G222gat & G426gat;
  assign new_G1197gat = G222gat & G443gat;
  assign new_G1200gat = G222gat & G460gat;
  assign new_G1203gat = G222gat & G477gat;
  assign new_G1206gat = G222gat & G494gat;
  assign new_G1209gat = G222gat & G511gat;
  assign new_G1212gat = G222gat & G528gat;
  assign new_G1215gat = G239gat & G273gat;
  assign new_G1218gat = G239gat & G290gat;
  assign new_G1221gat = G239gat & G307gat;
  assign new_G1224gat = G239gat & G324gat;
  assign new_G1227gat = G239gat & G341gat;
  assign new_G1230gat = G239gat & G358gat;
  assign new_G1233gat = G239gat & G375gat;
  assign new_G1236gat = G239gat & G392gat;
  assign new_G1239gat = G239gat & G409gat;
  assign new_G1242gat = G239gat & G426gat;
  assign new_G1245gat = G239gat & G443gat;
  assign new_G1248gat = G239gat & G460gat;
  assign new_G1251gat = G239gat & G477gat;
  assign new_G1254gat = G239gat & G494gat;
  assign new_G1257gat = G239gat & G511gat;
  assign new_G1260gat = G239gat & G528gat;
  assign new_G1263gat = G256gat & G273gat;
  assign new_G1266gat = G256gat & G290gat;
  assign new_G1269gat = G256gat & G307gat;
  assign new_G1272gat = G256gat & G324gat;
  assign new_G1275gat = G256gat & G341gat;
  assign new_G1278gat = G256gat & G358gat;
  assign new_G1281gat = G256gat & G375gat;
  assign new_G1284gat = G256gat & G392gat;
  assign new_G1287gat = G256gat & G409gat;
  assign new_G1290gat = G256gat & G426gat;
  assign new_G1293gat = G256gat & G443gat;
  assign new_G1296gat = G256gat & G460gat;
  assign new_G1299gat = G256gat & G477gat;
  assign new_G1302gat = G256gat & G494gat;
  assign new_G1305gat = G256gat & G511gat;
  assign new_G1308gat = G256gat & G528gat;
  assign new_G1311gat = ~new_G591gat;
  assign new_G1315gat = ~new_G639gat;
  assign new_G1319gat = ~new_G687gat;
  assign new_G1323gat = ~new_G735gat;
  assign new_G1327gat = ~new_G783gat;
  assign new_G1331gat = ~new_G831gat;
  assign new_G1335gat = ~new_G879gat;
  assign new_G1339gat = ~new_G927gat;
  assign new_G1343gat = ~new_G975gat;
  assign new_G1347gat = ~new_G1023gat;
  assign new_G1351gat = ~new_G1071gat;
  assign new_G1355gat = ~new_G1119gat;
  assign new_G1359gat = ~new_G1167gat;
  assign new_G1363gat = ~new_G1215gat;
  assign new_G1367gat = ~new_G1263gat;
  assign new_G1371gat = ~new_G591gat & ~new_G1311gat;
  assign new_G1372gat = ~new_G1311gat;
  assign new_G1373gat = ~new_G639gat & ~new_G1315gat;
  assign new_G1374gat = ~new_G1315gat;
  assign new_G1375gat = ~new_G687gat & ~new_G1319gat;
  assign new_G1376gat = ~new_G1319gat;
  assign new_G1377gat = ~new_G735gat & ~new_G1323gat;
  assign new_G1378gat = ~new_G1323gat;
  assign new_G1379gat = ~new_G783gat & ~new_G1327gat;
  assign new_G1380gat = ~new_G1327gat;
  assign new_G1381gat = ~new_G831gat & ~new_G1331gat;
  assign new_G1382gat = ~new_G1331gat;
  assign new_G1383gat = ~new_G879gat & ~new_G1335gat;
  assign new_G1384gat = ~new_G1335gat;
  assign new_G1385gat = ~new_G927gat & ~new_G1339gat;
  assign new_G1386gat = ~new_G1339gat;
  assign new_G1387gat = ~new_G975gat & ~new_G1343gat;
  assign new_G1388gat = ~new_G1343gat;
  assign new_G1389gat = ~new_G1023gat & ~new_G1347gat;
  assign new_G1390gat = ~new_G1347gat;
  assign new_G1391gat = ~new_G1071gat & ~new_G1351gat;
  assign new_G1392gat = ~new_G1351gat;
  assign new_G1393gat = ~new_G1119gat & ~new_G1355gat;
  assign new_G1394gat = ~new_G1355gat;
  assign new_G1395gat = ~new_G1167gat & ~new_G1359gat;
  assign new_G1396gat = ~new_G1359gat;
  assign new_G1397gat = ~new_G1215gat & ~new_G1363gat;
  assign new_G1398gat = ~new_G1363gat;
  assign new_G1399gat = ~new_G1263gat & ~new_G1367gat;
  assign new_G1400gat = ~new_G1367gat;
  assign new_G1401gat = ~new_G1371gat & ~new_G1372gat;
  assign new_G1404gat = ~new_G1373gat & ~new_G1374gat;
  assign new_G1407gat = ~new_G1375gat & ~new_G1376gat;
  assign new_G1410gat = ~new_G1377gat & ~new_G1378gat;
  assign new_G1413gat = ~new_G1379gat & ~new_G1380gat;
  assign new_G1416gat = ~new_G1381gat & ~new_G1382gat;
  assign new_G1419gat = ~new_G1383gat & ~new_G1384gat;
  assign new_G1422gat = ~new_G1385gat & ~new_G1386gat;
  assign new_G1425gat = ~new_G1387gat & ~new_G1388gat;
  assign new_G1428gat = ~new_G1389gat & ~new_G1390gat;
  assign new_G1431gat = ~new_G1391gat & ~new_G1392gat;
  assign new_G1434gat = ~new_G1393gat & ~new_G1394gat;
  assign new_G1437gat = ~new_G1395gat & ~new_G1396gat;
  assign new_G1440gat = ~new_G1397gat & ~new_G1398gat;
  assign new_G1443gat = ~new_G1399gat & ~new_G1400gat;
  assign new_G1446gat = ~new_G1401gat & ~new_G546gat;
  assign new_G1450gat = ~new_G1404gat & ~new_G594gat;
  assign new_G1454gat = ~new_G1407gat & ~new_G642gat;
  assign new_G1458gat = ~new_G1410gat & ~new_G690gat;
  assign new_G1462gat = ~new_G1413gat & ~new_G738gat;
  assign new_G1466gat = ~new_G1416gat & ~new_G786gat;
  assign new_G1470gat = ~new_G1419gat & ~new_G834gat;
  assign new_G1474gat = ~new_G1422gat & ~new_G882gat;
  assign new_G1478gat = ~new_G1425gat & ~new_G930gat;
  assign new_G1482gat = ~new_G1428gat & ~new_G978gat;
  assign new_G1486gat = ~new_G1431gat & ~new_G1026gat;
  assign new_G1490gat = ~new_G1434gat & ~new_G1074gat;
  assign new_G1494gat = ~new_G1437gat & ~new_G1122gat;
  assign new_G1498gat = ~new_G1440gat & ~new_G1170gat;
  assign new_G1502gat = ~new_G1443gat & ~new_G1218gat;
  assign new_G1506gat = ~new_G1401gat & ~new_G1446gat;
  assign new_G1507gat = ~new_G1446gat & ~new_G546gat;
  assign new_G1508gat = ~new_G1311gat & ~new_G1446gat;
  assign new_G1511gat = ~new_G1404gat & ~new_G1450gat;
  assign new_G1512gat = ~new_G1450gat & ~new_G594gat;
  assign new_G1513gat = ~new_G1315gat & ~new_G1450gat;
  assign new_G1516gat = ~new_G1407gat & ~new_G1454gat;
  assign new_G1517gat = ~new_G1454gat & ~new_G642gat;
  assign new_G1518gat = ~new_G1319gat & ~new_G1454gat;
  assign new_G1521gat = ~new_G1410gat & ~new_G1458gat;
  assign new_G1522gat = ~new_G1458gat & ~new_G690gat;
  assign new_G1523gat = ~new_G1323gat & ~new_G1458gat;
  assign new_G1526gat = ~new_G1413gat & ~new_G1462gat;
  assign new_G1527gat = ~new_G1462gat & ~new_G738gat;
  assign new_G1528gat = ~new_G1327gat & ~new_G1462gat;
  assign new_G1531gat = ~new_G1416gat & ~new_G1466gat;
  assign new_G1532gat = ~new_G1466gat & ~new_G786gat;
  assign new_G1533gat = ~new_G1331gat & ~new_G1466gat;
  assign new_G1536gat = ~new_G1419gat & ~new_G1470gat;
  assign new_G1537gat = ~new_G1470gat & ~new_G834gat;
  assign new_G1538gat = ~new_G1335gat & ~new_G1470gat;
  assign new_G1541gat = ~new_G1422gat & ~new_G1474gat;
  assign new_G1542gat = ~new_G1474gat & ~new_G882gat;
  assign new_G1543gat = ~new_G1339gat & ~new_G1474gat;
  assign new_G1546gat = ~new_G1425gat & ~new_G1478gat;
  assign new_G1547gat = ~new_G1478gat & ~new_G930gat;
  assign new_G1548gat = ~new_G1343gat & ~new_G1478gat;
  assign new_G1551gat = ~new_G1428gat & ~new_G1482gat;
  assign new_G1552gat = ~new_G1482gat & ~new_G978gat;
  assign new_G1553gat = ~new_G1347gat & ~new_G1482gat;
  assign new_G1556gat = ~new_G1431gat & ~new_G1486gat;
  assign new_G1557gat = ~new_G1486gat & ~new_G1026gat;
  assign new_G1558gat = ~new_G1351gat & ~new_G1486gat;
  assign new_G1561gat = ~new_G1434gat & ~new_G1490gat;
  assign new_G1562gat = ~new_G1490gat & ~new_G1074gat;
  assign new_G1563gat = ~new_G1355gat & ~new_G1490gat;
  assign new_G1566gat = ~new_G1437gat & ~new_G1494gat;
  assign new_G1567gat = ~new_G1494gat & ~new_G1122gat;
  assign new_G1568gat = ~new_G1359gat & ~new_G1494gat;
  assign new_G1571gat = ~new_G1440gat & ~new_G1498gat;
  assign new_G1572gat = ~new_G1498gat & ~new_G1170gat;
  assign new_G1573gat = ~new_G1363gat & ~new_G1498gat;
  assign new_G1576gat = ~new_G1443gat & ~new_G1502gat;
  assign new_G1577gat = ~new_G1502gat & ~new_G1218gat;
  assign new_G1578gat = ~new_G1367gat & ~new_G1502gat;
  assign G1581gat = ~new_G1506gat & ~new_G1507gat;
  assign new_G1582gat = ~new_G1511gat & ~new_G1512gat;
  assign new_G1585gat = ~new_G1516gat & ~new_G1517gat;
  assign new_G1588gat = ~new_G1521gat & ~new_G1522gat;
  assign new_G1591gat = ~new_G1526gat & ~new_G1527gat;
  assign new_G1594gat = ~new_G1531gat & ~new_G1532gat;
  assign new_G1597gat = ~new_G1536gat & ~new_G1537gat;
  assign new_G1600gat = ~new_G1541gat & ~new_G1542gat;
  assign new_G1603gat = ~new_G1546gat & ~new_G1547gat;
  assign new_G1606gat = ~new_G1551gat & ~new_G1552gat;
  assign new_G1609gat = ~new_G1556gat & ~new_G1557gat;
  assign new_G1612gat = ~new_G1561gat & ~new_G1562gat;
  assign new_G1615gat = ~new_G1566gat & ~new_G1567gat;
  assign new_G1618gat = ~new_G1571gat & ~new_G1572gat;
  assign new_G1621gat = ~new_G1576gat & ~new_G1577gat;
  assign new_G1624gat = ~new_G1266gat & ~new_G1578gat;
  assign new_G1628gat = ~new_G1582gat & ~new_G1508gat;
  assign new_G1632gat = ~new_G1585gat & ~new_G1513gat;
  assign new_G1636gat = ~new_G1588gat & ~new_G1518gat;
  assign new_G1640gat = ~new_G1591gat & ~new_G1523gat;
  assign new_G1644gat = ~new_G1594gat & ~new_G1528gat;
  assign new_G1648gat = ~new_G1597gat & ~new_G1533gat;
  assign new_G1652gat = ~new_G1600gat & ~new_G1538gat;
  assign new_G1656gat = ~new_G1603gat & ~new_G1543gat;
  assign new_G1660gat = ~new_G1606gat & ~new_G1548gat;
  assign new_G1664gat = ~new_G1609gat & ~new_G1553gat;
  assign new_G1668gat = ~new_G1612gat & ~new_G1558gat;
  assign new_G1672gat = ~new_G1615gat & ~new_G1563gat;
  assign new_G1676gat = ~new_G1618gat & ~new_G1568gat;
  assign new_G1680gat = ~new_G1621gat & ~new_G1573gat;
  assign new_G1684gat = ~new_G1266gat & ~new_G1624gat;
  assign new_G1685gat = ~new_G1624gat & ~new_G1578gat;
  assign new_G1686gat = ~new_G1582gat & ~new_G1628gat;
  assign new_G1687gat = ~new_G1628gat & ~new_G1508gat;
  assign new_G1688gat = ~new_G1585gat & ~new_G1632gat;
  assign new_G1689gat = ~new_G1632gat & ~new_G1513gat;
  assign new_G1690gat = ~new_G1588gat & ~new_G1636gat;
  assign new_G1691gat = ~new_G1636gat & ~new_G1518gat;
  assign new_G1692gat = ~new_G1591gat & ~new_G1640gat;
  assign new_G1693gat = ~new_G1640gat & ~new_G1523gat;
  assign new_G1694gat = ~new_G1594gat & ~new_G1644gat;
  assign new_G1695gat = ~new_G1644gat & ~new_G1528gat;
  assign new_G1696gat = ~new_G1597gat & ~new_G1648gat;
  assign new_G1697gat = ~new_G1648gat & ~new_G1533gat;
  assign new_G1698gat = ~new_G1600gat & ~new_G1652gat;
  assign new_G1699gat = ~new_G1652gat & ~new_G1538gat;
  assign new_G1700gat = ~new_G1603gat & ~new_G1656gat;
  assign new_G1701gat = ~new_G1656gat & ~new_G1543gat;
  assign new_G1702gat = ~new_G1606gat & ~new_G1660gat;
  assign new_G1703gat = ~new_G1660gat & ~new_G1548gat;
  assign new_G1704gat = ~new_G1609gat & ~new_G1664gat;
  assign new_G1705gat = ~new_G1664gat & ~new_G1553gat;
  assign new_G1706gat = ~new_G1612gat & ~new_G1668gat;
  assign new_G1707gat = ~new_G1668gat & ~new_G1558gat;
  assign new_G1708gat = ~new_G1615gat & ~new_G1672gat;
  assign new_G1709gat = ~new_G1672gat & ~new_G1563gat;
  assign new_G1710gat = ~new_G1618gat & ~new_G1676gat;
  assign new_G1711gat = ~new_G1676gat & ~new_G1568gat;
  assign new_G1712gat = ~new_G1621gat & ~new_G1680gat;
  assign new_G1713gat = ~new_G1680gat & ~new_G1573gat;
  assign new_G1714gat = ~new_G1684gat & ~new_G1685gat;
  assign new_G1717gat = ~new_G1686gat & ~new_G1687gat;
  assign new_G1720gat = ~new_G1688gat & ~new_G1689gat;
  assign new_G1723gat = ~new_G1690gat & ~new_G1691gat;
  assign new_G1726gat = ~new_G1692gat & ~new_G1693gat;
  assign new_G1729gat = ~new_G1694gat & ~new_G1695gat;
  assign new_G1732gat = ~new_G1696gat & ~new_G1697gat;
  assign new_G1735gat = ~new_G1698gat & ~new_G1699gat;
  assign new_G1738gat = ~new_G1700gat & ~new_G1701gat;
  assign new_G1741gat = ~new_G1702gat & ~new_G1703gat;
  assign new_G1744gat = ~new_G1704gat & ~new_G1705gat;
  assign new_G1747gat = ~new_G1706gat & ~new_G1707gat;
  assign new_G1750gat = ~new_G1708gat & ~new_G1709gat;
  assign new_G1753gat = ~new_G1710gat & ~new_G1711gat;
  assign new_G1756gat = ~new_G1712gat & ~new_G1713gat;
  assign new_G1759gat = ~new_G1714gat & ~new_G1221gat;
  assign new_G1763gat = ~new_G1717gat & ~new_G549gat;
  assign new_G1767gat = ~new_G1720gat & ~new_G597gat;
  assign new_G1771gat = ~new_G1723gat & ~new_G645gat;
  assign new_G1775gat = ~new_G1726gat & ~new_G693gat;
  assign new_G1779gat = ~new_G1729gat & ~new_G741gat;
  assign new_G1783gat = ~new_G1732gat & ~new_G789gat;
  assign new_G1787gat = ~new_G1735gat & ~new_G837gat;
  assign new_G1791gat = ~new_G1738gat & ~new_G885gat;
  assign new_G1795gat = ~new_G1741gat & ~new_G933gat;
  assign new_G1799gat = ~new_G1744gat & ~new_G981gat;
  assign new_G1803gat = ~new_G1747gat & ~new_G1029gat;
  assign new_G1807gat = ~new_G1750gat & ~new_G1077gat;
  assign new_G1811gat = ~new_G1753gat & ~new_G1125gat;
  assign new_G1815gat = ~new_G1756gat & ~new_G1173gat;
  assign new_G1819gat = ~new_G1714gat & ~new_G1759gat;
  assign new_G1820gat = ~new_G1759gat & ~new_G1221gat;
  assign new_G1821gat = ~new_G1624gat & ~new_G1759gat;
  assign new_G1824gat = ~new_G1717gat & ~new_G1763gat;
  assign new_G1825gat = ~new_G1763gat & ~new_G549gat;
  assign new_G1826gat = ~new_G1628gat & ~new_G1763gat;
  assign new_G1829gat = ~new_G1720gat & ~new_G1767gat;
  assign new_G1830gat = ~new_G1767gat & ~new_G597gat;
  assign new_G1831gat = ~new_G1632gat & ~new_G1767gat;
  assign new_G1834gat = ~new_G1723gat & ~new_G1771gat;
  assign new_G1835gat = ~new_G1771gat & ~new_G645gat;
  assign new_G1836gat = ~new_G1636gat & ~new_G1771gat;
  assign new_G1839gat = ~new_G1726gat & ~new_G1775gat;
  assign new_G1840gat = ~new_G1775gat & ~new_G693gat;
  assign new_G1841gat = ~new_G1640gat & ~new_G1775gat;
  assign new_G1844gat = ~new_G1729gat & ~new_G1779gat;
  assign new_G1845gat = ~new_G1779gat & ~new_G741gat;
  assign new_G1846gat = ~new_G1644gat & ~new_G1779gat;
  assign new_G1849gat = ~new_G1732gat & ~new_G1783gat;
  assign new_G1850gat = ~new_G1783gat & ~new_G789gat;
  assign new_G1851gat = ~new_G1648gat & ~new_G1783gat;
  assign new_G1854gat = ~new_G1735gat & ~new_G1787gat;
  assign new_G1855gat = ~new_G1787gat & ~new_G837gat;
  assign new_G1856gat = ~new_G1652gat & ~new_G1787gat;
  assign new_G1859gat = ~new_G1738gat & ~new_G1791gat;
  assign new_G1860gat = ~new_G1791gat & ~new_G885gat;
  assign new_G1861gat = ~new_G1656gat & ~new_G1791gat;
  assign new_G1864gat = ~new_G1741gat & ~new_G1795gat;
  assign new_G1865gat = ~new_G1795gat & ~new_G933gat;
  assign new_G1866gat = ~new_G1660gat & ~new_G1795gat;
  assign new_G1869gat = ~new_G1744gat & ~new_G1799gat;
  assign new_G1870gat = ~new_G1799gat & ~new_G981gat;
  assign new_G1871gat = ~new_G1664gat & ~new_G1799gat;
  assign new_G1874gat = ~new_G1747gat & ~new_G1803gat;
  assign new_G1875gat = ~new_G1803gat & ~new_G1029gat;
  assign new_G1876gat = ~new_G1668gat & ~new_G1803gat;
  assign new_G1879gat = ~new_G1750gat & ~new_G1807gat;
  assign new_G1880gat = ~new_G1807gat & ~new_G1077gat;
  assign new_G1881gat = ~new_G1672gat & ~new_G1807gat;
  assign new_G1884gat = ~new_G1753gat & ~new_G1811gat;
  assign new_G1885gat = ~new_G1811gat & ~new_G1125gat;
  assign new_G1886gat = ~new_G1676gat & ~new_G1811gat;
  assign new_G1889gat = ~new_G1756gat & ~new_G1815gat;
  assign new_G1890gat = ~new_G1815gat & ~new_G1173gat;
  assign new_G1891gat = ~new_G1680gat & ~new_G1815gat;
  assign new_G1894gat = ~new_G1819gat & ~new_G1820gat;
  assign new_G1897gat = ~new_G1269gat & ~new_G1821gat;
  assign G1901gat = ~new_G1824gat & ~new_G1825gat;
  assign new_G1902gat = ~new_G1829gat & ~new_G1830gat;
  assign new_G1905gat = ~new_G1834gat & ~new_G1835gat;
  assign new_G1908gat = ~new_G1839gat & ~new_G1840gat;
  assign new_G1911gat = ~new_G1844gat & ~new_G1845gat;
  assign new_G1914gat = ~new_G1849gat & ~new_G1850gat;
  assign new_G1917gat = ~new_G1854gat & ~new_G1855gat;
  assign new_G1920gat = ~new_G1859gat & ~new_G1860gat;
  assign new_G1923gat = ~new_G1864gat & ~new_G1865gat;
  assign new_G1926gat = ~new_G1869gat & ~new_G1870gat;
  assign new_G1929gat = ~new_G1874gat & ~new_G1875gat;
  assign new_G1932gat = ~new_G1879gat & ~new_G1880gat;
  assign new_G1935gat = ~new_G1884gat & ~new_G1885gat;
  assign new_G1938gat = ~new_G1889gat & ~new_G1890gat;
  assign new_G1941gat = ~new_G1894gat & ~new_G1891gat;
  assign new_G1945gat = ~new_G1269gat & ~new_G1897gat;
  assign new_G1946gat = ~new_G1897gat & ~new_G1821gat;
  assign new_G1947gat = ~new_G1902gat & ~new_G1826gat;
  assign new_G1951gat = ~new_G1905gat & ~new_G1831gat;
  assign new_G1955gat = ~new_G1908gat & ~new_G1836gat;
  assign new_G1959gat = ~new_G1911gat & ~new_G1841gat;
  assign new_G1963gat = ~new_G1914gat & ~new_G1846gat;
  assign new_G1967gat = ~new_G1917gat & ~new_G1851gat;
  assign new_G1971gat = ~new_G1920gat & ~new_G1856gat;
  assign new_G1975gat = ~new_G1923gat & ~new_G1861gat;
  assign new_G1979gat = ~new_G1926gat & ~new_G1866gat;
  assign new_G1983gat = ~new_G1929gat & ~new_G1871gat;
  assign new_G1987gat = ~new_G1932gat & ~new_G1876gat;
  assign new_G1991gat = ~new_G1935gat & ~new_G1881gat;
  assign new_G1995gat = ~new_G1938gat & ~new_G1886gat;
  assign new_G1999gat = ~new_G1894gat & ~new_G1941gat;
  assign new_G2000gat = ~new_G1941gat & ~new_G1891gat;
  assign new_G2001gat = ~new_G1945gat & ~new_G1946gat;
  assign new_G2004gat = ~new_G1902gat & ~new_G1947gat;
  assign new_G2005gat = ~new_G1947gat & ~new_G1826gat;
  assign new_G2006gat = ~new_G1905gat & ~new_G1951gat;
  assign new_G2007gat = ~new_G1951gat & ~new_G1831gat;
  assign new_G2008gat = ~new_G1908gat & ~new_G1955gat;
  assign new_G2009gat = ~new_G1955gat & ~new_G1836gat;
  assign new_G2010gat = ~new_G1911gat & ~new_G1959gat;
  assign new_G2011gat = ~new_G1959gat & ~new_G1841gat;
  assign new_G2012gat = ~new_G1914gat & ~new_G1963gat;
  assign new_G2013gat = ~new_G1963gat & ~new_G1846gat;
  assign new_G2014gat = ~new_G1917gat & ~new_G1967gat;
  assign new_G2015gat = ~new_G1967gat & ~new_G1851gat;
  assign new_G2016gat = ~new_G1920gat & ~new_G1971gat;
  assign new_G2017gat = ~new_G1971gat & ~new_G1856gat;
  assign new_G2018gat = ~new_G1923gat & ~new_G1975gat;
  assign new_G2019gat = ~new_G1975gat & ~new_G1861gat;
  assign new_G2020gat = ~new_G1926gat & ~new_G1979gat;
  assign new_G2021gat = ~new_G1979gat & ~new_G1866gat;
  assign new_G2022gat = ~new_G1929gat & ~new_G1983gat;
  assign new_G2023gat = ~new_G1983gat & ~new_G1871gat;
  assign new_G2024gat = ~new_G1932gat & ~new_G1987gat;
  assign new_G2025gat = ~new_G1987gat & ~new_G1876gat;
  assign new_G2026gat = ~new_G1935gat & ~new_G1991gat;
  assign new_G2027gat = ~new_G1991gat & ~new_G1881gat;
  assign new_G2028gat = ~new_G1938gat & ~new_G1995gat;
  assign new_G2029gat = ~new_G1995gat & ~new_G1886gat;
  assign new_G2030gat = ~new_G1999gat & ~new_G2000gat;
  assign new_G2033gat = ~new_G2001gat & ~new_G1224gat;
  assign new_G2037gat = ~new_G2004gat & ~new_G2005gat;
  assign new_G2040gat = ~new_G2006gat & ~new_G2007gat;
  assign new_G2043gat = ~new_G2008gat & ~new_G2009gat;
  assign new_G2046gat = ~new_G2010gat & ~new_G2011gat;
  assign new_G2049gat = ~new_G2012gat & ~new_G2013gat;
  assign new_G2052gat = ~new_G2014gat & ~new_G2015gat;
  assign new_G2055gat = ~new_G2016gat & ~new_G2017gat;
  assign new_G2058gat = ~new_G2018gat & ~new_G2019gat;
  assign new_G2061gat = ~new_G2020gat & ~new_G2021gat;
  assign new_G2064gat = ~new_G2022gat & ~new_G2023gat;
  assign new_G2067gat = ~new_G2024gat & ~new_G2025gat;
  assign new_G2070gat = ~new_G2026gat & ~new_G2027gat;
  assign new_G2073gat = ~new_G2028gat & ~new_G2029gat;
  assign new_G2076gat = ~new_G2030gat & ~new_G1176gat;
  assign new_G2080gat = ~new_G2001gat & ~new_G2033gat;
  assign new_G2081gat = ~new_G2033gat & ~new_G1224gat;
  assign new_G2082gat = ~new_G1897gat & ~new_G2033gat;
  assign new_G2085gat = ~new_G2037gat & ~new_G552gat;
  assign new_G2089gat = ~new_G2040gat & ~new_G600gat;
  assign new_G2093gat = ~new_G2043gat & ~new_G648gat;
  assign new_G2097gat = ~new_G2046gat & ~new_G696gat;
  assign new_G2101gat = ~new_G2049gat & ~new_G744gat;
  assign new_G2105gat = ~new_G2052gat & ~new_G792gat;
  assign new_G2109gat = ~new_G2055gat & ~new_G840gat;
  assign new_G2113gat = ~new_G2058gat & ~new_G888gat;
  assign new_G2117gat = ~new_G2061gat & ~new_G936gat;
  assign new_G2121gat = ~new_G2064gat & ~new_G984gat;
  assign new_G2125gat = ~new_G2067gat & ~new_G1032gat;
  assign new_G2129gat = ~new_G2070gat & ~new_G1080gat;
  assign new_G2133gat = ~new_G2073gat & ~new_G1128gat;
  assign new_G2137gat = ~new_G2030gat & ~new_G2076gat;
  assign new_G2138gat = ~new_G2076gat & ~new_G1176gat;
  assign new_G2139gat = ~new_G1941gat & ~new_G2076gat;
  assign new_G2142gat = ~new_G2080gat & ~new_G2081gat;
  assign new_G2145gat = ~new_G1272gat & ~new_G2082gat;
  assign new_G2149gat = ~new_G2037gat & ~new_G2085gat;
  assign new_G2150gat = ~new_G2085gat & ~new_G552gat;
  assign new_G2151gat = ~new_G1947gat & ~new_G2085gat;
  assign new_G2154gat = ~new_G2040gat & ~new_G2089gat;
  assign new_G2155gat = ~new_G2089gat & ~new_G600gat;
  assign new_G2156gat = ~new_G1951gat & ~new_G2089gat;
  assign new_G2159gat = ~new_G2043gat & ~new_G2093gat;
  assign new_G2160gat = ~new_G2093gat & ~new_G648gat;
  assign new_G2161gat = ~new_G1955gat & ~new_G2093gat;
  assign new_G2164gat = ~new_G2046gat & ~new_G2097gat;
  assign new_G2165gat = ~new_G2097gat & ~new_G696gat;
  assign new_G2166gat = ~new_G1959gat & ~new_G2097gat;
  assign new_G2169gat = ~new_G2049gat & ~new_G2101gat;
  assign new_G2170gat = ~new_G2101gat & ~new_G744gat;
  assign new_G2171gat = ~new_G1963gat & ~new_G2101gat;
  assign new_G2174gat = ~new_G2052gat & ~new_G2105gat;
  assign new_G2175gat = ~new_G2105gat & ~new_G792gat;
  assign new_G2176gat = ~new_G1967gat & ~new_G2105gat;
  assign new_G2179gat = ~new_G2055gat & ~new_G2109gat;
  assign new_G2180gat = ~new_G2109gat & ~new_G840gat;
  assign new_G2181gat = ~new_G1971gat & ~new_G2109gat;
  assign new_G2184gat = ~new_G2058gat & ~new_G2113gat;
  assign new_G2185gat = ~new_G2113gat & ~new_G888gat;
  assign new_G2186gat = ~new_G1975gat & ~new_G2113gat;
  assign new_G2189gat = ~new_G2061gat & ~new_G2117gat;
  assign new_G2190gat = ~new_G2117gat & ~new_G936gat;
  assign new_G2191gat = ~new_G1979gat & ~new_G2117gat;
  assign new_G2194gat = ~new_G2064gat & ~new_G2121gat;
  assign new_G2195gat = ~new_G2121gat & ~new_G984gat;
  assign new_G2196gat = ~new_G1983gat & ~new_G2121gat;
  assign new_G2199gat = ~new_G2067gat & ~new_G2125gat;
  assign new_G2200gat = ~new_G2125gat & ~new_G1032gat;
  assign new_G2201gat = ~new_G1987gat & ~new_G2125gat;
  assign new_G2204gat = ~new_G2070gat & ~new_G2129gat;
  assign new_G2205gat = ~new_G2129gat & ~new_G1080gat;
  assign new_G2206gat = ~new_G1991gat & ~new_G2129gat;
  assign new_G2209gat = ~new_G2073gat & ~new_G2133gat;
  assign new_G2210gat = ~new_G2133gat & ~new_G1128gat;
  assign new_G2211gat = ~new_G1995gat & ~new_G2133gat;
  assign new_G2214gat = ~new_G2137gat & ~new_G2138gat;
  assign new_G2217gat = ~new_G2142gat & ~new_G2139gat;
  assign new_G2221gat = ~new_G1272gat & ~new_G2145gat;
  assign new_G2222gat = ~new_G2145gat & ~new_G2082gat;
  assign G2223gat = ~new_G2149gat & ~new_G2150gat;
  assign new_G2224gat = ~new_G2154gat & ~new_G2155gat;
  assign new_G2227gat = ~new_G2159gat & ~new_G2160gat;
  assign new_G2230gat = ~new_G2164gat & ~new_G2165gat;
  assign new_G2233gat = ~new_G2169gat & ~new_G2170gat;
  assign new_G2236gat = ~new_G2174gat & ~new_G2175gat;
  assign new_G2239gat = ~new_G2179gat & ~new_G2180gat;
  assign new_G2242gat = ~new_G2184gat & ~new_G2185gat;
  assign new_G2245gat = ~new_G2189gat & ~new_G2190gat;
  assign new_G2248gat = ~new_G2194gat & ~new_G2195gat;
  assign new_G2251gat = ~new_G2199gat & ~new_G2200gat;
  assign new_G2254gat = ~new_G2204gat & ~new_G2205gat;
  assign new_G2257gat = ~new_G2209gat & ~new_G2210gat;
  assign new_G2260gat = ~new_G2214gat & ~new_G2211gat;
  assign new_G2264gat = ~new_G2142gat & ~new_G2217gat;
  assign new_G2265gat = ~new_G2217gat & ~new_G2139gat;
  assign new_G2266gat = ~new_G2221gat & ~new_G2222gat;
  assign new_G2269gat = ~new_G2224gat & ~new_G2151gat;
  assign new_G2273gat = ~new_G2227gat & ~new_G2156gat;
  assign new_G2277gat = ~new_G2230gat & ~new_G2161gat;
  assign new_G2281gat = ~new_G2233gat & ~new_G2166gat;
  assign new_G2285gat = ~new_G2236gat & ~new_G2171gat;
  assign new_G2289gat = ~new_G2239gat & ~new_G2176gat;
  assign new_G2293gat = ~new_G2242gat & ~new_G2181gat;
  assign new_G2297gat = ~new_G2245gat & ~new_G2186gat;
  assign new_G2301gat = ~new_G2248gat & ~new_G2191gat;
  assign new_G2305gat = ~new_G2251gat & ~new_G2196gat;
  assign new_G2309gat = ~new_G2254gat & ~new_G2201gat;
  assign new_G2313gat = ~new_G2257gat & ~new_G2206gat;
  assign new_G2317gat = ~new_G2214gat & ~new_G2260gat;
  assign new_G2318gat = ~new_G2260gat & ~new_G2211gat;
  assign new_G2319gat = ~new_G2264gat & ~new_G2265gat;
  assign new_G2322gat = ~new_G2266gat & ~new_G1227gat;
  assign new_G2326gat = ~new_G2224gat & ~new_G2269gat;
  assign new_G2327gat = ~new_G2269gat & ~new_G2151gat;
  assign new_G2328gat = ~new_G2227gat & ~new_G2273gat;
  assign new_G2329gat = ~new_G2273gat & ~new_G2156gat;
  assign new_G2330gat = ~new_G2230gat & ~new_G2277gat;
  assign new_G2331gat = ~new_G2277gat & ~new_G2161gat;
  assign new_G2332gat = ~new_G2233gat & ~new_G2281gat;
  assign new_G2333gat = ~new_G2281gat & ~new_G2166gat;
  assign new_G2334gat = ~new_G2236gat & ~new_G2285gat;
  assign new_G2335gat = ~new_G2285gat & ~new_G2171gat;
  assign new_G2336gat = ~new_G2239gat & ~new_G2289gat;
  assign new_G2337gat = ~new_G2289gat & ~new_G2176gat;
  assign new_G2338gat = ~new_G2242gat & ~new_G2293gat;
  assign new_G2339gat = ~new_G2293gat & ~new_G2181gat;
  assign new_G2340gat = ~new_G2245gat & ~new_G2297gat;
  assign new_G2341gat = ~new_G2297gat & ~new_G2186gat;
  assign new_G2342gat = ~new_G2248gat & ~new_G2301gat;
  assign new_G2343gat = ~new_G2301gat & ~new_G2191gat;
  assign new_G2344gat = ~new_G2251gat & ~new_G2305gat;
  assign new_G2345gat = ~new_G2305gat & ~new_G2196gat;
  assign new_G2346gat = ~new_G2254gat & ~new_G2309gat;
  assign new_G2347gat = ~new_G2309gat & ~new_G2201gat;
  assign new_G2348gat = ~new_G2257gat & ~new_G2313gat;
  assign new_G2349gat = ~new_G2313gat & ~new_G2206gat;
  assign new_G2350gat = ~new_G2317gat & ~new_G2318gat;
  assign new_G2353gat = ~new_G2319gat & ~new_G1179gat;
  assign new_G2357gat = ~new_G2266gat & ~new_G2322gat;
  assign new_G2358gat = ~new_G2322gat & ~new_G1227gat;
  assign new_G2359gat = ~new_G2145gat & ~new_G2322gat;
  assign new_G2362gat = ~new_G2326gat & ~new_G2327gat;
  assign new_G2365gat = ~new_G2328gat & ~new_G2329gat;
  assign new_G2368gat = ~new_G2330gat & ~new_G2331gat;
  assign new_G2371gat = ~new_G2332gat & ~new_G2333gat;
  assign new_G2374gat = ~new_G2334gat & ~new_G2335gat;
  assign new_G2377gat = ~new_G2336gat & ~new_G2337gat;
  assign new_G2380gat = ~new_G2338gat & ~new_G2339gat;
  assign new_G2383gat = ~new_G2340gat & ~new_G2341gat;
  assign new_G2386gat = ~new_G2342gat & ~new_G2343gat;
  assign new_G2389gat = ~new_G2344gat & ~new_G2345gat;
  assign new_G2392gat = ~new_G2346gat & ~new_G2347gat;
  assign new_G2395gat = ~new_G2348gat & ~new_G2349gat;
  assign new_G2398gat = ~new_G2350gat & ~new_G1131gat;
  assign new_G2402gat = ~new_G2319gat & ~new_G2353gat;
  assign new_G2403gat = ~new_G2353gat & ~new_G1179gat;
  assign new_G2404gat = ~new_G2217gat & ~new_G2353gat;
  assign new_G2407gat = ~new_G2357gat & ~new_G2358gat;
  assign new_G2410gat = ~new_G1275gat & ~new_G2359gat;
  assign new_G2414gat = ~new_G2362gat & ~new_G555gat;
  assign new_G2418gat = ~new_G2365gat & ~new_G603gat;
  assign new_G2422gat = ~new_G2368gat & ~new_G651gat;
  assign new_G2426gat = ~new_G2371gat & ~new_G699gat;
  assign new_G2430gat = ~new_G2374gat & ~new_G747gat;
  assign new_G2434gat = ~new_G2377gat & ~new_G795gat;
  assign new_G2438gat = ~new_G2380gat & ~new_G843gat;
  assign new_G2442gat = ~new_G2383gat & ~new_G891gat;
  assign new_G2446gat = ~new_G2386gat & ~new_G939gat;
  assign new_G2450gat = ~new_G2389gat & ~new_G987gat;
  assign new_G2454gat = ~new_G2392gat & ~new_G1035gat;
  assign new_G2458gat = ~new_G2395gat & ~new_G1083gat;
  assign new_G2462gat = ~new_G2350gat & ~new_G2398gat;
  assign new_G2463gat = ~new_G2398gat & ~new_G1131gat;
  assign new_G2464gat = ~new_G2260gat & ~new_G2398gat;
  assign new_G2467gat = ~new_G2402gat & ~new_G2403gat;
  assign new_G2470gat = ~new_G2407gat & ~new_G2404gat;
  assign new_G2474gat = ~new_G1275gat & ~new_G2410gat;
  assign new_G2475gat = ~new_G2410gat & ~new_G2359gat;
  assign new_G2476gat = ~new_G2362gat & ~new_G2414gat;
  assign new_G2477gat = ~new_G2414gat & ~new_G555gat;
  assign new_G2478gat = ~new_G2269gat & ~new_G2414gat;
  assign new_G2481gat = ~new_G2365gat & ~new_G2418gat;
  assign new_G2482gat = ~new_G2418gat & ~new_G603gat;
  assign new_G2483gat = ~new_G2273gat & ~new_G2418gat;
  assign new_G2486gat = ~new_G2368gat & ~new_G2422gat;
  assign new_G2487gat = ~new_G2422gat & ~new_G651gat;
  assign new_G2488gat = ~new_G2277gat & ~new_G2422gat;
  assign new_G2491gat = ~new_G2371gat & ~new_G2426gat;
  assign new_G2492gat = ~new_G2426gat & ~new_G699gat;
  assign new_G2493gat = ~new_G2281gat & ~new_G2426gat;
  assign new_G2496gat = ~new_G2374gat & ~new_G2430gat;
  assign new_G2497gat = ~new_G2430gat & ~new_G747gat;
  assign new_G2498gat = ~new_G2285gat & ~new_G2430gat;
  assign new_G2501gat = ~new_G2377gat & ~new_G2434gat;
  assign new_G2502gat = ~new_G2434gat & ~new_G795gat;
  assign new_G2503gat = ~new_G2289gat & ~new_G2434gat;
  assign new_G2506gat = ~new_G2380gat & ~new_G2438gat;
  assign new_G2507gat = ~new_G2438gat & ~new_G843gat;
  assign new_G2508gat = ~new_G2293gat & ~new_G2438gat;
  assign new_G2511gat = ~new_G2383gat & ~new_G2442gat;
  assign new_G2512gat = ~new_G2442gat & ~new_G891gat;
  assign new_G2513gat = ~new_G2297gat & ~new_G2442gat;
  assign new_G2516gat = ~new_G2386gat & ~new_G2446gat;
  assign new_G2517gat = ~new_G2446gat & ~new_G939gat;
  assign new_G2518gat = ~new_G2301gat & ~new_G2446gat;
  assign new_G2521gat = ~new_G2389gat & ~new_G2450gat;
  assign new_G2522gat = ~new_G2450gat & ~new_G987gat;
  assign new_G2523gat = ~new_G2305gat & ~new_G2450gat;
  assign new_G2526gat = ~new_G2392gat & ~new_G2454gat;
  assign new_G2527gat = ~new_G2454gat & ~new_G1035gat;
  assign new_G2528gat = ~new_G2309gat & ~new_G2454gat;
  assign new_G2531gat = ~new_G2395gat & ~new_G2458gat;
  assign new_G2532gat = ~new_G2458gat & ~new_G1083gat;
  assign new_G2533gat = ~new_G2313gat & ~new_G2458gat;
  assign new_G2536gat = ~new_G2462gat & ~new_G2463gat;
  assign new_G2539gat = ~new_G2467gat & ~new_G2464gat;
  assign new_G2543gat = ~new_G2407gat & ~new_G2470gat;
  assign new_G2544gat = ~new_G2470gat & ~new_G2404gat;
  assign new_G2545gat = ~new_G2474gat & ~new_G2475gat;
  assign G2548gat = ~new_G2476gat & ~new_G2477gat;
  assign new_G2549gat = ~new_G2481gat & ~new_G2482gat;
  assign new_G2552gat = ~new_G2486gat & ~new_G2487gat;
  assign new_G2555gat = ~new_G2491gat & ~new_G2492gat;
  assign new_G2558gat = ~new_G2496gat & ~new_G2497gat;
  assign new_G2561gat = ~new_G2501gat & ~new_G2502gat;
  assign new_G2564gat = ~new_G2506gat & ~new_G2507gat;
  assign new_G2567gat = ~new_G2511gat & ~new_G2512gat;
  assign new_G2570gat = ~new_G2516gat & ~new_G2517gat;
  assign new_G2573gat = ~new_G2521gat & ~new_G2522gat;
  assign new_G2576gat = ~new_G2526gat & ~new_G2527gat;
  assign new_G2579gat = ~new_G2531gat & ~new_G2532gat;
  assign new_G2582gat = ~new_G2536gat & ~new_G2533gat;
  assign new_G2586gat = ~new_G2467gat & ~new_G2539gat;
  assign new_G2587gat = ~new_G2539gat & ~new_G2464gat;
  assign new_G2588gat = ~new_G2543gat & ~new_G2544gat;
  assign new_G2591gat = ~new_G2545gat & ~new_G1230gat;
  assign new_G2595gat = ~new_G2549gat & ~new_G2478gat;
  assign new_G2599gat = ~new_G2552gat & ~new_G2483gat;
  assign new_G2603gat = ~new_G2555gat & ~new_G2488gat;
  assign new_G2607gat = ~new_G2558gat & ~new_G2493gat;
  assign new_G2611gat = ~new_G2561gat & ~new_G2498gat;
  assign new_G2615gat = ~new_G2564gat & ~new_G2503gat;
  assign new_G2619gat = ~new_G2567gat & ~new_G2508gat;
  assign new_G2623gat = ~new_G2570gat & ~new_G2513gat;
  assign new_G2627gat = ~new_G2573gat & ~new_G2518gat;
  assign new_G2631gat = ~new_G2576gat & ~new_G2523gat;
  assign new_G2635gat = ~new_G2579gat & ~new_G2528gat;
  assign new_G2639gat = ~new_G2536gat & ~new_G2582gat;
  assign new_G2640gat = ~new_G2582gat & ~new_G2533gat;
  assign new_G2641gat = ~new_G2586gat & ~new_G2587gat;
  assign new_G2644gat = ~new_G2588gat & ~new_G1182gat;
  assign new_G2648gat = ~new_G2545gat & ~new_G2591gat;
  assign new_G2649gat = ~new_G2591gat & ~new_G1230gat;
  assign new_G2650gat = ~new_G2410gat & ~new_G2591gat;
  assign new_G2653gat = ~new_G2549gat & ~new_G2595gat;
  assign new_G2654gat = ~new_G2595gat & ~new_G2478gat;
  assign new_G2655gat = ~new_G2552gat & ~new_G2599gat;
  assign new_G2656gat = ~new_G2599gat & ~new_G2483gat;
  assign new_G2657gat = ~new_G2555gat & ~new_G2603gat;
  assign new_G2658gat = ~new_G2603gat & ~new_G2488gat;
  assign new_G2659gat = ~new_G2558gat & ~new_G2607gat;
  assign new_G2660gat = ~new_G2607gat & ~new_G2493gat;
  assign new_G2661gat = ~new_G2561gat & ~new_G2611gat;
  assign new_G2662gat = ~new_G2611gat & ~new_G2498gat;
  assign new_G2663gat = ~new_G2564gat & ~new_G2615gat;
  assign new_G2664gat = ~new_G2615gat & ~new_G2503gat;
  assign new_G2665gat = ~new_G2567gat & ~new_G2619gat;
  assign new_G2666gat = ~new_G2619gat & ~new_G2508gat;
  assign new_G2667gat = ~new_G2570gat & ~new_G2623gat;
  assign new_G2668gat = ~new_G2623gat & ~new_G2513gat;
  assign new_G2669gat = ~new_G2573gat & ~new_G2627gat;
  assign new_G2670gat = ~new_G2627gat & ~new_G2518gat;
  assign new_G2671gat = ~new_G2576gat & ~new_G2631gat;
  assign new_G2672gat = ~new_G2631gat & ~new_G2523gat;
  assign new_G2673gat = ~new_G2579gat & ~new_G2635gat;
  assign new_G2674gat = ~new_G2635gat & ~new_G2528gat;
  assign new_G2675gat = ~new_G2639gat & ~new_G2640gat;
  assign new_G2678gat = ~new_G2641gat & ~new_G1134gat;
  assign new_G2682gat = ~new_G2588gat & ~new_G2644gat;
  assign new_G2683gat = ~new_G2644gat & ~new_G1182gat;
  assign new_G2684gat = ~new_G2470gat & ~new_G2644gat;
  assign new_G2687gat = ~new_G2648gat & ~new_G2649gat;
  assign new_G2690gat = ~new_G1278gat & ~new_G2650gat;
  assign new_G2694gat = ~new_G2653gat & ~new_G2654gat;
  assign new_G2697gat = ~new_G2655gat & ~new_G2656gat;
  assign new_G2700gat = ~new_G2657gat & ~new_G2658gat;
  assign new_G2703gat = ~new_G2659gat & ~new_G2660gat;
  assign new_G2706gat = ~new_G2661gat & ~new_G2662gat;
  assign new_G2709gat = ~new_G2663gat & ~new_G2664gat;
  assign new_G2712gat = ~new_G2665gat & ~new_G2666gat;
  assign new_G2715gat = ~new_G2667gat & ~new_G2668gat;
  assign new_G2718gat = ~new_G2669gat & ~new_G2670gat;
  assign new_G2721gat = ~new_G2671gat & ~new_G2672gat;
  assign new_G2724gat = ~new_G2673gat & ~new_G2674gat;
  assign new_G2727gat = ~new_G2675gat & ~new_G1086gat;
  assign new_G2731gat = ~new_G2641gat & ~new_G2678gat;
  assign new_G2732gat = ~new_G2678gat & ~new_G1134gat;
  assign new_G2733gat = ~new_G2539gat & ~new_G2678gat;
  assign new_G2736gat = ~new_G2682gat & ~new_G2683gat;
  assign new_G2739gat = ~new_G2687gat & ~new_G2684gat;
  assign new_G2743gat = ~new_G1278gat & ~new_G2690gat;
  assign new_G2744gat = ~new_G2690gat & ~new_G2650gat;
  assign new_G2745gat = ~new_G2694gat & ~new_G558gat;
  assign new_G2749gat = ~new_G2697gat & ~new_G606gat;
  assign new_G2753gat = ~new_G2700gat & ~new_G654gat;
  assign new_G2757gat = ~new_G2703gat & ~new_G702gat;
  assign new_G2761gat = ~new_G2706gat & ~new_G750gat;
  assign new_G2765gat = ~new_G2709gat & ~new_G798gat;
  assign new_G2769gat = ~new_G2712gat & ~new_G846gat;
  assign new_G2773gat = ~new_G2715gat & ~new_G894gat;
  assign new_G2777gat = ~new_G2718gat & ~new_G942gat;
  assign new_G2781gat = ~new_G2721gat & ~new_G990gat;
  assign new_G2785gat = ~new_G2724gat & ~new_G1038gat;
  assign new_G2789gat = ~new_G2675gat & ~new_G2727gat;
  assign new_G2790gat = ~new_G2727gat & ~new_G1086gat;
  assign new_G2791gat = ~new_G2582gat & ~new_G2727gat;
  assign new_G2794gat = ~new_G2731gat & ~new_G2732gat;
  assign new_G2797gat = ~new_G2736gat & ~new_G2733gat;
  assign new_G2801gat = ~new_G2687gat & ~new_G2739gat;
  assign new_G2802gat = ~new_G2739gat & ~new_G2684gat;
  assign new_G2803gat = ~new_G2743gat & ~new_G2744gat;
  assign new_G2806gat = ~new_G2694gat & ~new_G2745gat;
  assign new_G2807gat = ~new_G2745gat & ~new_G558gat;
  assign new_G2808gat = ~new_G2595gat & ~new_G2745gat;
  assign new_G2811gat = ~new_G2697gat & ~new_G2749gat;
  assign new_G2812gat = ~new_G2749gat & ~new_G606gat;
  assign new_G2813gat = ~new_G2599gat & ~new_G2749gat;
  assign new_G2816gat = ~new_G2700gat & ~new_G2753gat;
  assign new_G2817gat = ~new_G2753gat & ~new_G654gat;
  assign new_G2818gat = ~new_G2603gat & ~new_G2753gat;
  assign new_G2821gat = ~new_G2703gat & ~new_G2757gat;
  assign new_G2822gat = ~new_G2757gat & ~new_G702gat;
  assign new_G2823gat = ~new_G2607gat & ~new_G2757gat;
  assign new_G2826gat = ~new_G2706gat & ~new_G2761gat;
  assign new_G2827gat = ~new_G2761gat & ~new_G750gat;
  assign new_G2828gat = ~new_G2611gat & ~new_G2761gat;
  assign new_G2831gat = ~new_G2709gat & ~new_G2765gat;
  assign new_G2832gat = ~new_G2765gat & ~new_G798gat;
  assign new_G2833gat = ~new_G2615gat & ~new_G2765gat;
  assign new_G2836gat = ~new_G2712gat & ~new_G2769gat;
  assign new_G2837gat = ~new_G2769gat & ~new_G846gat;
  assign new_G2838gat = ~new_G2619gat & ~new_G2769gat;
  assign new_G2841gat = ~new_G2715gat & ~new_G2773gat;
  assign new_G2842gat = ~new_G2773gat & ~new_G894gat;
  assign new_G2843gat = ~new_G2623gat & ~new_G2773gat;
  assign new_G2846gat = ~new_G2718gat & ~new_G2777gat;
  assign new_G2847gat = ~new_G2777gat & ~new_G942gat;
  assign new_G2848gat = ~new_G2627gat & ~new_G2777gat;
  assign new_G2851gat = ~new_G2721gat & ~new_G2781gat;
  assign new_G2852gat = ~new_G2781gat & ~new_G990gat;
  assign new_G2853gat = ~new_G2631gat & ~new_G2781gat;
  assign new_G2856gat = ~new_G2724gat & ~new_G2785gat;
  assign new_G2857gat = ~new_G2785gat & ~new_G1038gat;
  assign new_G2858gat = ~new_G2635gat & ~new_G2785gat;
  assign new_G2861gat = ~new_G2789gat & ~new_G2790gat;
  assign new_G2864gat = ~new_G2794gat & ~new_G2791gat;
  assign new_G2868gat = ~new_G2736gat & ~new_G2797gat;
  assign new_G2869gat = ~new_G2797gat & ~new_G2733gat;
  assign new_G2870gat = ~new_G2801gat & ~new_G2802gat;
  assign new_G2873gat = ~new_G2803gat & ~new_G1233gat;
  assign G2877gat = ~new_G2806gat & ~new_G2807gat;
  assign new_G2878gat = ~new_G2811gat & ~new_G2812gat;
  assign new_G2881gat = ~new_G2816gat & ~new_G2817gat;
  assign new_G2884gat = ~new_G2821gat & ~new_G2822gat;
  assign new_G2887gat = ~new_G2826gat & ~new_G2827gat;
  assign new_G2890gat = ~new_G2831gat & ~new_G2832gat;
  assign new_G2893gat = ~new_G2836gat & ~new_G2837gat;
  assign new_G2896gat = ~new_G2841gat & ~new_G2842gat;
  assign new_G2899gat = ~new_G2846gat & ~new_G2847gat;
  assign new_G2902gat = ~new_G2851gat & ~new_G2852gat;
  assign new_G2905gat = ~new_G2856gat & ~new_G2857gat;
  assign new_G2908gat = ~new_G2861gat & ~new_G2858gat;
  assign new_G2912gat = ~new_G2794gat & ~new_G2864gat;
  assign new_G2913gat = ~new_G2864gat & ~new_G2791gat;
  assign new_G2914gat = ~new_G2868gat & ~new_G2869gat;
  assign new_G2917gat = ~new_G2870gat & ~new_G1185gat;
  assign new_G2921gat = ~new_G2803gat & ~new_G2873gat;
  assign new_G2922gat = ~new_G2873gat & ~new_G1233gat;
  assign new_G2923gat = ~new_G2690gat & ~new_G2873gat;
  assign new_G2926gat = ~new_G2878gat & ~new_G2808gat;
  assign new_G2930gat = ~new_G2881gat & ~new_G2813gat;
  assign new_G2934gat = ~new_G2884gat & ~new_G2818gat;
  assign new_G2938gat = ~new_G2887gat & ~new_G2823gat;
  assign new_G2942gat = ~new_G2890gat & ~new_G2828gat;
  assign new_G2946gat = ~new_G2893gat & ~new_G2833gat;
  assign new_G2950gat = ~new_G2896gat & ~new_G2838gat;
  assign new_G2954gat = ~new_G2899gat & ~new_G2843gat;
  assign new_G2958gat = ~new_G2902gat & ~new_G2848gat;
  assign new_G2962gat = ~new_G2905gat & ~new_G2853gat;
  assign new_G2966gat = ~new_G2861gat & ~new_G2908gat;
  assign new_G2967gat = ~new_G2908gat & ~new_G2858gat;
  assign new_G2968gat = ~new_G2912gat & ~new_G2913gat;
  assign new_G2971gat = ~new_G2914gat & ~new_G1137gat;
  assign new_G2975gat = ~new_G2870gat & ~new_G2917gat;
  assign new_G2976gat = ~new_G2917gat & ~new_G1185gat;
  assign new_G2977gat = ~new_G2739gat & ~new_G2917gat;
  assign new_G2980gat = ~new_G2921gat & ~new_G2922gat;
  assign new_G2983gat = ~new_G1281gat & ~new_G2923gat;
  assign new_G2987gat = ~new_G2878gat & ~new_G2926gat;
  assign new_G2988gat = ~new_G2926gat & ~new_G2808gat;
  assign new_G2989gat = ~new_G2881gat & ~new_G2930gat;
  assign new_G2990gat = ~new_G2930gat & ~new_G2813gat;
  assign new_G2991gat = ~new_G2884gat & ~new_G2934gat;
  assign new_G2992gat = ~new_G2934gat & ~new_G2818gat;
  assign new_G2993gat = ~new_G2887gat & ~new_G2938gat;
  assign new_G2994gat = ~new_G2938gat & ~new_G2823gat;
  assign new_G2995gat = ~new_G2890gat & ~new_G2942gat;
  assign new_G2996gat = ~new_G2942gat & ~new_G2828gat;
  assign new_G2997gat = ~new_G2893gat & ~new_G2946gat;
  assign new_G2998gat = ~new_G2946gat & ~new_G2833gat;
  assign new_G2999gat = ~new_G2896gat & ~new_G2950gat;
  assign new_G3000gat = ~new_G2950gat & ~new_G2838gat;
  assign new_G3001gat = ~new_G2899gat & ~new_G2954gat;
  assign new_G3002gat = ~new_G2954gat & ~new_G2843gat;
  assign new_G3003gat = ~new_G2902gat & ~new_G2958gat;
  assign new_G3004gat = ~new_G2958gat & ~new_G2848gat;
  assign new_G3005gat = ~new_G2905gat & ~new_G2962gat;
  assign new_G3006gat = ~new_G2962gat & ~new_G2853gat;
  assign new_G3007gat = ~new_G2966gat & ~new_G2967gat;
  assign new_G3010gat = ~new_G2968gat & ~new_G1089gat;
  assign new_G3014gat = ~new_G2914gat & ~new_G2971gat;
  assign new_G3015gat = ~new_G2971gat & ~new_G1137gat;
  assign new_G3016gat = ~new_G2797gat & ~new_G2971gat;
  assign new_G3019gat = ~new_G2975gat & ~new_G2976gat;
  assign new_G3022gat = ~new_G2980gat & ~new_G2977gat;
  assign new_G3026gat = ~new_G1281gat & ~new_G2983gat;
  assign new_G3027gat = ~new_G2983gat & ~new_G2923gat;
  assign new_G3028gat = ~new_G2987gat & ~new_G2988gat;
  assign new_G3031gat = ~new_G2989gat & ~new_G2990gat;
  assign new_G3034gat = ~new_G2991gat & ~new_G2992gat;
  assign new_G3037gat = ~new_G2993gat & ~new_G2994gat;
  assign new_G3040gat = ~new_G2995gat & ~new_G2996gat;
  assign new_G3043gat = ~new_G2997gat & ~new_G2998gat;
  assign new_G3046gat = ~new_G2999gat & ~new_G3000gat;
  assign new_G3049gat = ~new_G3001gat & ~new_G3002gat;
  assign new_G3052gat = ~new_G3003gat & ~new_G3004gat;
  assign new_G3055gat = ~new_G3005gat & ~new_G3006gat;
  assign new_G3058gat = ~new_G3007gat & ~new_G1041gat;
  assign new_G3062gat = ~new_G2968gat & ~new_G3010gat;
  assign new_G3063gat = ~new_G3010gat & ~new_G1089gat;
  assign new_G3064gat = ~new_G2864gat & ~new_G3010gat;
  assign new_G3067gat = ~new_G3014gat & ~new_G3015gat;
  assign new_G3070gat = ~new_G3019gat & ~new_G3016gat;
  assign new_G3074gat = ~new_G2980gat & ~new_G3022gat;
  assign new_G3075gat = ~new_G3022gat & ~new_G2977gat;
  assign new_G3076gat = ~new_G3026gat & ~new_G3027gat;
  assign new_G3079gat = ~new_G3028gat & ~new_G561gat;
  assign new_G3083gat = ~new_G3031gat & ~new_G609gat;
  assign new_G3087gat = ~new_G3034gat & ~new_G657gat;
  assign new_G3091gat = ~new_G3037gat & ~new_G705gat;
  assign new_G3095gat = ~new_G3040gat & ~new_G753gat;
  assign new_G3099gat = ~new_G3043gat & ~new_G801gat;
  assign new_G3103gat = ~new_G3046gat & ~new_G849gat;
  assign new_G3107gat = ~new_G3049gat & ~new_G897gat;
  assign new_G3111gat = ~new_G3052gat & ~new_G945gat;
  assign new_G3115gat = ~new_G3055gat & ~new_G993gat;
  assign new_G3119gat = ~new_G3007gat & ~new_G3058gat;
  assign new_G3120gat = ~new_G3058gat & ~new_G1041gat;
  assign new_G3121gat = ~new_G2908gat & ~new_G3058gat;
  assign new_G3124gat = ~new_G3062gat & ~new_G3063gat;
  assign new_G3127gat = ~new_G3067gat & ~new_G3064gat;
  assign new_G3131gat = ~new_G3019gat & ~new_G3070gat;
  assign new_G3132gat = ~new_G3070gat & ~new_G3016gat;
  assign new_G3133gat = ~new_G3074gat & ~new_G3075gat;
  assign new_G3136gat = ~new_G3076gat & ~new_G1236gat;
  assign new_G3140gat = ~new_G3028gat & ~new_G3079gat;
  assign new_G3141gat = ~new_G3079gat & ~new_G561gat;
  assign new_G3142gat = ~new_G2926gat & ~new_G3079gat;
  assign new_G3145gat = ~new_G3031gat & ~new_G3083gat;
  assign new_G3146gat = ~new_G3083gat & ~new_G609gat;
  assign new_G3147gat = ~new_G2930gat & ~new_G3083gat;
  assign new_G3150gat = ~new_G3034gat & ~new_G3087gat;
  assign new_G3151gat = ~new_G3087gat & ~new_G657gat;
  assign new_G3152gat = ~new_G2934gat & ~new_G3087gat;
  assign new_G3155gat = ~new_G3037gat & ~new_G3091gat;
  assign new_G3156gat = ~new_G3091gat & ~new_G705gat;
  assign new_G3157gat = ~new_G2938gat & ~new_G3091gat;
  assign new_G3160gat = ~new_G3040gat & ~new_G3095gat;
  assign new_G3161gat = ~new_G3095gat & ~new_G753gat;
  assign new_G3162gat = ~new_G2942gat & ~new_G3095gat;
  assign new_G3165gat = ~new_G3043gat & ~new_G3099gat;
  assign new_G3166gat = ~new_G3099gat & ~new_G801gat;
  assign new_G3167gat = ~new_G2946gat & ~new_G3099gat;
  assign new_G3170gat = ~new_G3046gat & ~new_G3103gat;
  assign new_G3171gat = ~new_G3103gat & ~new_G849gat;
  assign new_G3172gat = ~new_G2950gat & ~new_G3103gat;
  assign new_G3175gat = ~new_G3049gat & ~new_G3107gat;
  assign new_G3176gat = ~new_G3107gat & ~new_G897gat;
  assign new_G3177gat = ~new_G2954gat & ~new_G3107gat;
  assign new_G3180gat = ~new_G3052gat & ~new_G3111gat;
  assign new_G3181gat = ~new_G3111gat & ~new_G945gat;
  assign new_G3182gat = ~new_G2958gat & ~new_G3111gat;
  assign new_G3185gat = ~new_G3055gat & ~new_G3115gat;
  assign new_G3186gat = ~new_G3115gat & ~new_G993gat;
  assign new_G3187gat = ~new_G2962gat & ~new_G3115gat;
  assign new_G3190gat = ~new_G3119gat & ~new_G3120gat;
  assign new_G3193gat = ~new_G3124gat & ~new_G3121gat;
  assign new_G3197gat = ~new_G3067gat & ~new_G3127gat;
  assign new_G3198gat = ~new_G3127gat & ~new_G3064gat;
  assign new_G3199gat = ~new_G3131gat & ~new_G3132gat;
  assign new_G3202gat = ~new_G3133gat & ~new_G1188gat;
  assign new_G3206gat = ~new_G3076gat & ~new_G3136gat;
  assign new_G3207gat = ~new_G3136gat & ~new_G1236gat;
  assign new_G3208gat = ~new_G2983gat & ~new_G3136gat;
  assign G3211gat = ~new_G3140gat & ~new_G3141gat;
  assign new_G3212gat = ~new_G3145gat & ~new_G3146gat;
  assign new_G3215gat = ~new_G3150gat & ~new_G3151gat;
  assign new_G3218gat = ~new_G3155gat & ~new_G3156gat;
  assign new_G3221gat = ~new_G3160gat & ~new_G3161gat;
  assign new_G3224gat = ~new_G3165gat & ~new_G3166gat;
  assign new_G3227gat = ~new_G3170gat & ~new_G3171gat;
  assign new_G3230gat = ~new_G3175gat & ~new_G3176gat;
  assign new_G3233gat = ~new_G3180gat & ~new_G3181gat;
  assign new_G3236gat = ~new_G3185gat & ~new_G3186gat;
  assign new_G3239gat = ~new_G3190gat & ~new_G3187gat;
  assign new_G3243gat = ~new_G3124gat & ~new_G3193gat;
  assign new_G3244gat = ~new_G3193gat & ~new_G3121gat;
  assign new_G3245gat = ~new_G3197gat & ~new_G3198gat;
  assign new_G3248gat = ~new_G3199gat & ~new_G1140gat;
  assign new_G3252gat = ~new_G3133gat & ~new_G3202gat;
  assign new_G3253gat = ~new_G3202gat & ~new_G1188gat;
  assign new_G3254gat = ~new_G3022gat & ~new_G3202gat;
  assign new_G3257gat = ~new_G3206gat & ~new_G3207gat;
  assign new_G3260gat = ~new_G1284gat & ~new_G3208gat;
  assign new_G3264gat = ~new_G3212gat & ~new_G3142gat;
  assign new_G3268gat = ~new_G3215gat & ~new_G3147gat;
  assign new_G3272gat = ~new_G3218gat & ~new_G3152gat;
  assign new_G3276gat = ~new_G3221gat & ~new_G3157gat;
  assign new_G3280gat = ~new_G3224gat & ~new_G3162gat;
  assign new_G3284gat = ~new_G3227gat & ~new_G3167gat;
  assign new_G3288gat = ~new_G3230gat & ~new_G3172gat;
  assign new_G3292gat = ~new_G3233gat & ~new_G3177gat;
  assign new_G3296gat = ~new_G3236gat & ~new_G3182gat;
  assign new_G3300gat = ~new_G3190gat & ~new_G3239gat;
  assign new_G3301gat = ~new_G3239gat & ~new_G3187gat;
  assign new_G3302gat = ~new_G3243gat & ~new_G3244gat;
  assign new_G3305gat = ~new_G3245gat & ~new_G1092gat;
  assign new_G3309gat = ~new_G3199gat & ~new_G3248gat;
  assign new_G3310gat = ~new_G3248gat & ~new_G1140gat;
  assign new_G3311gat = ~new_G3070gat & ~new_G3248gat;
  assign new_G3314gat = ~new_G3252gat & ~new_G3253gat;
  assign new_G3317gat = ~new_G3257gat & ~new_G3254gat;
  assign new_G3321gat = ~new_G1284gat & ~new_G3260gat;
  assign new_G3322gat = ~new_G3260gat & ~new_G3208gat;
  assign new_G3323gat = ~new_G3212gat & ~new_G3264gat;
  assign new_G3324gat = ~new_G3264gat & ~new_G3142gat;
  assign new_G3325gat = ~new_G3215gat & ~new_G3268gat;
  assign new_G3326gat = ~new_G3268gat & ~new_G3147gat;
  assign new_G3327gat = ~new_G3218gat & ~new_G3272gat;
  assign new_G3328gat = ~new_G3272gat & ~new_G3152gat;
  assign new_G3329gat = ~new_G3221gat & ~new_G3276gat;
  assign new_G3330gat = ~new_G3276gat & ~new_G3157gat;
  assign new_G3331gat = ~new_G3224gat & ~new_G3280gat;
  assign new_G3332gat = ~new_G3280gat & ~new_G3162gat;
  assign new_G3333gat = ~new_G3227gat & ~new_G3284gat;
  assign new_G3334gat = ~new_G3284gat & ~new_G3167gat;
  assign new_G3335gat = ~new_G3230gat & ~new_G3288gat;
  assign new_G3336gat = ~new_G3288gat & ~new_G3172gat;
  assign new_G3337gat = ~new_G3233gat & ~new_G3292gat;
  assign new_G3338gat = ~new_G3292gat & ~new_G3177gat;
  assign new_G3339gat = ~new_G3236gat & ~new_G3296gat;
  assign new_G3340gat = ~new_G3296gat & ~new_G3182gat;
  assign new_G3341gat = ~new_G3300gat & ~new_G3301gat;
  assign new_G3344gat = ~new_G3302gat & ~new_G1044gat;
  assign new_G3348gat = ~new_G3245gat & ~new_G3305gat;
  assign new_G3349gat = ~new_G3305gat & ~new_G1092gat;
  assign new_G3350gat = ~new_G3127gat & ~new_G3305gat;
  assign new_G3353gat = ~new_G3309gat & ~new_G3310gat;
  assign new_G3356gat = ~new_G3314gat & ~new_G3311gat;
  assign new_G3360gat = ~new_G3257gat & ~new_G3317gat;
  assign new_G3361gat = ~new_G3317gat & ~new_G3254gat;
  assign new_G3362gat = ~new_G3321gat & ~new_G3322gat;
  assign new_G3365gat = ~new_G3323gat & ~new_G3324gat;
  assign new_G3368gat = ~new_G3325gat & ~new_G3326gat;
  assign new_G3371gat = ~new_G3327gat & ~new_G3328gat;
  assign new_G3374gat = ~new_G3329gat & ~new_G3330gat;
  assign new_G3377gat = ~new_G3331gat & ~new_G3332gat;
  assign new_G3380gat = ~new_G3333gat & ~new_G3334gat;
  assign new_G3383gat = ~new_G3335gat & ~new_G3336gat;
  assign new_G3386gat = ~new_G3337gat & ~new_G3338gat;
  assign new_G3389gat = ~new_G3339gat & ~new_G3340gat;
  assign new_G3392gat = ~new_G3341gat & ~new_G996gat;
  assign new_G3396gat = ~new_G3302gat & ~new_G3344gat;
  assign new_G3397gat = ~new_G3344gat & ~new_G1044gat;
  assign new_G3398gat = ~new_G3193gat & ~new_G3344gat;
  assign new_G3401gat = ~new_G3348gat & ~new_G3349gat;
  assign new_G3404gat = ~new_G3353gat & ~new_G3350gat;
  assign new_G3408gat = ~new_G3314gat & ~new_G3356gat;
  assign new_G3409gat = ~new_G3356gat & ~new_G3311gat;
  assign new_G3410gat = ~new_G3360gat & ~new_G3361gat;
  assign new_G3413gat = ~new_G3362gat & ~new_G1239gat;
  assign new_G3417gat = ~new_G3365gat & ~new_G564gat;
  assign new_G3421gat = ~new_G3368gat & ~new_G612gat;
  assign new_G3425gat = ~new_G3371gat & ~new_G660gat;
  assign new_G3429gat = ~new_G3374gat & ~new_G708gat;
  assign new_G3433gat = ~new_G3377gat & ~new_G756gat;
  assign new_G3437gat = ~new_G3380gat & ~new_G804gat;
  assign new_G3441gat = ~new_G3383gat & ~new_G852gat;
  assign new_G3445gat = ~new_G3386gat & ~new_G900gat;
  assign new_G3449gat = ~new_G3389gat & ~new_G948gat;
  assign new_G3453gat = ~new_G3341gat & ~new_G3392gat;
  assign new_G3454gat = ~new_G3392gat & ~new_G996gat;
  assign new_G3455gat = ~new_G3239gat & ~new_G3392gat;
  assign new_G3458gat = ~new_G3396gat & ~new_G3397gat;
  assign new_G3461gat = ~new_G3401gat & ~new_G3398gat;
  assign new_G3465gat = ~new_G3353gat & ~new_G3404gat;
  assign new_G3466gat = ~new_G3404gat & ~new_G3350gat;
  assign new_G3467gat = ~new_G3408gat & ~new_G3409gat;
  assign new_G3470gat = ~new_G3410gat & ~new_G1191gat;
  assign new_G3474gat = ~new_G3362gat & ~new_G3413gat;
  assign new_G3475gat = ~new_G3413gat & ~new_G1239gat;
  assign new_G3476gat = ~new_G3260gat & ~new_G3413gat;
  assign new_G3479gat = ~new_G3365gat & ~new_G3417gat;
  assign new_G3480gat = ~new_G3417gat & ~new_G564gat;
  assign new_G3481gat = ~new_G3264gat & ~new_G3417gat;
  assign new_G3484gat = ~new_G3368gat & ~new_G3421gat;
  assign new_G3485gat = ~new_G3421gat & ~new_G612gat;
  assign new_G3486gat = ~new_G3268gat & ~new_G3421gat;
  assign new_G3489gat = ~new_G3371gat & ~new_G3425gat;
  assign new_G3490gat = ~new_G3425gat & ~new_G660gat;
  assign new_G3491gat = ~new_G3272gat & ~new_G3425gat;
  assign new_G3494gat = ~new_G3374gat & ~new_G3429gat;
  assign new_G3495gat = ~new_G3429gat & ~new_G708gat;
  assign new_G3496gat = ~new_G3276gat & ~new_G3429gat;
  assign new_G3499gat = ~new_G3377gat & ~new_G3433gat;
  assign new_G3500gat = ~new_G3433gat & ~new_G756gat;
  assign new_G3501gat = ~new_G3280gat & ~new_G3433gat;
  assign new_G3504gat = ~new_G3380gat & ~new_G3437gat;
  assign new_G3505gat = ~new_G3437gat & ~new_G804gat;
  assign new_G3506gat = ~new_G3284gat & ~new_G3437gat;
  assign new_G3509gat = ~new_G3383gat & ~new_G3441gat;
  assign new_G3510gat = ~new_G3441gat & ~new_G852gat;
  assign new_G3511gat = ~new_G3288gat & ~new_G3441gat;
  assign new_G3514gat = ~new_G3386gat & ~new_G3445gat;
  assign new_G3515gat = ~new_G3445gat & ~new_G900gat;
  assign new_G3516gat = ~new_G3292gat & ~new_G3445gat;
  assign new_G3519gat = ~new_G3389gat & ~new_G3449gat;
  assign new_G3520gat = ~new_G3449gat & ~new_G948gat;
  assign new_G3521gat = ~new_G3296gat & ~new_G3449gat;
  assign new_G3524gat = ~new_G3453gat & ~new_G3454gat;
  assign new_G3527gat = ~new_G3458gat & ~new_G3455gat;
  assign new_G3531gat = ~new_G3401gat & ~new_G3461gat;
  assign new_G3532gat = ~new_G3461gat & ~new_G3398gat;
  assign new_G3533gat = ~new_G3465gat & ~new_G3466gat;
  assign new_G3536gat = ~new_G3467gat & ~new_G1143gat;
  assign new_G3540gat = ~new_G3410gat & ~new_G3470gat;
  assign new_G3541gat = ~new_G3470gat & ~new_G1191gat;
  assign new_G3542gat = ~new_G3317gat & ~new_G3470gat;
  assign new_G3545gat = ~new_G3474gat & ~new_G3475gat;
  assign new_G3548gat = ~new_G1287gat & ~new_G3476gat;
  assign G3552gat = ~new_G3479gat & ~new_G3480gat;
  assign new_G3553gat = ~new_G3484gat & ~new_G3485gat;
  assign new_G3556gat = ~new_G3489gat & ~new_G3490gat;
  assign new_G3559gat = ~new_G3494gat & ~new_G3495gat;
  assign new_G3562gat = ~new_G3499gat & ~new_G3500gat;
  assign new_G3565gat = ~new_G3504gat & ~new_G3505gat;
  assign new_G3568gat = ~new_G3509gat & ~new_G3510gat;
  assign new_G3571gat = ~new_G3514gat & ~new_G3515gat;
  assign new_G3574gat = ~new_G3519gat & ~new_G3520gat;
  assign new_G3577gat = ~new_G3524gat & ~new_G3521gat;
  assign new_G3581gat = ~new_G3458gat & ~new_G3527gat;
  assign new_G3582gat = ~new_G3527gat & ~new_G3455gat;
  assign new_G3583gat = ~new_G3531gat & ~new_G3532gat;
  assign new_G3586gat = ~new_G3533gat & ~new_G1095gat;
  assign new_G3590gat = ~new_G3467gat & ~new_G3536gat;
  assign new_G3591gat = ~new_G3536gat & ~new_G1143gat;
  assign new_G3592gat = ~new_G3356gat & ~new_G3536gat;
  assign new_G3595gat = ~new_G3540gat & ~new_G3541gat;
  assign new_G3598gat = ~new_G3545gat & ~new_G3542gat;
  assign new_G3602gat = ~new_G1287gat & ~new_G3548gat;
  assign new_G3603gat = ~new_G3548gat & ~new_G3476gat;
  assign new_G3604gat = ~new_G3553gat & ~new_G3481gat;
  assign new_G3608gat = ~new_G3556gat & ~new_G3486gat;
  assign new_G3612gat = ~new_G3559gat & ~new_G3491gat;
  assign new_G3616gat = ~new_G3562gat & ~new_G3496gat;
  assign new_G3620gat = ~new_G3565gat & ~new_G3501gat;
  assign new_G3624gat = ~new_G3568gat & ~new_G3506gat;
  assign new_G3628gat = ~new_G3571gat & ~new_G3511gat;
  assign new_G3632gat = ~new_G3574gat & ~new_G3516gat;
  assign new_G3636gat = ~new_G3524gat & ~new_G3577gat;
  assign new_G3637gat = ~new_G3577gat & ~new_G3521gat;
  assign new_G3638gat = ~new_G3581gat & ~new_G3582gat;
  assign new_G3641gat = ~new_G3583gat & ~new_G1047gat;
  assign new_G3645gat = ~new_G3533gat & ~new_G3586gat;
  assign new_G3646gat = ~new_G3586gat & ~new_G1095gat;
  assign new_G3647gat = ~new_G3404gat & ~new_G3586gat;
  assign new_G3650gat = ~new_G3590gat & ~new_G3591gat;
  assign new_G3653gat = ~new_G3595gat & ~new_G3592gat;
  assign new_G3657gat = ~new_G3545gat & ~new_G3598gat;
  assign new_G3658gat = ~new_G3598gat & ~new_G3542gat;
  assign new_G3659gat = ~new_G3602gat & ~new_G3603gat;
  assign new_G3662gat = ~new_G3553gat & ~new_G3604gat;
  assign new_G3663gat = ~new_G3604gat & ~new_G3481gat;
  assign new_G3664gat = ~new_G3556gat & ~new_G3608gat;
  assign new_G3665gat = ~new_G3608gat & ~new_G3486gat;
  assign new_G3666gat = ~new_G3559gat & ~new_G3612gat;
  assign new_G3667gat = ~new_G3612gat & ~new_G3491gat;
  assign new_G3668gat = ~new_G3562gat & ~new_G3616gat;
  assign new_G3669gat = ~new_G3616gat & ~new_G3496gat;
  assign new_G3670gat = ~new_G3565gat & ~new_G3620gat;
  assign new_G3671gat = ~new_G3620gat & ~new_G3501gat;
  assign new_G3672gat = ~new_G3568gat & ~new_G3624gat;
  assign new_G3673gat = ~new_G3624gat & ~new_G3506gat;
  assign new_G3674gat = ~new_G3571gat & ~new_G3628gat;
  assign new_G3675gat = ~new_G3628gat & ~new_G3511gat;
  assign new_G3676gat = ~new_G3574gat & ~new_G3632gat;
  assign new_G3677gat = ~new_G3632gat & ~new_G3516gat;
  assign new_G3678gat = ~new_G3636gat & ~new_G3637gat;
  assign new_G3681gat = ~new_G3638gat & ~new_G999gat;
  assign new_G3685gat = ~new_G3583gat & ~new_G3641gat;
  assign new_G3686gat = ~new_G3641gat & ~new_G1047gat;
  assign new_G3687gat = ~new_G3461gat & ~new_G3641gat;
  assign new_G3690gat = ~new_G3645gat & ~new_G3646gat;
  assign new_G3693gat = ~new_G3650gat & ~new_G3647gat;
  assign new_G3697gat = ~new_G3595gat & ~new_G3653gat;
  assign new_G3698gat = ~new_G3653gat & ~new_G3592gat;
  assign new_G3699gat = ~new_G3657gat & ~new_G3658gat;
  assign new_G3702gat = ~new_G3659gat & ~new_G1242gat;
  assign new_G3706gat = ~new_G3662gat & ~new_G3663gat;
  assign new_G3709gat = ~new_G3664gat & ~new_G3665gat;
  assign new_G3712gat = ~new_G3666gat & ~new_G3667gat;
  assign new_G3715gat = ~new_G3668gat & ~new_G3669gat;
  assign new_G3718gat = ~new_G3670gat & ~new_G3671gat;
  assign new_G3721gat = ~new_G3672gat & ~new_G3673gat;
  assign new_G3724gat = ~new_G3674gat & ~new_G3675gat;
  assign new_G3727gat = ~new_G3676gat & ~new_G3677gat;
  assign new_G3730gat = ~new_G3678gat & ~new_G951gat;
  assign new_G3734gat = ~new_G3638gat & ~new_G3681gat;
  assign new_G3735gat = ~new_G3681gat & ~new_G999gat;
  assign new_G3736gat = ~new_G3527gat & ~new_G3681gat;
  assign new_G3739gat = ~new_G3685gat & ~new_G3686gat;
  assign new_G3742gat = ~new_G3690gat & ~new_G3687gat;
  assign new_G3746gat = ~new_G3650gat & ~new_G3693gat;
  assign new_G3747gat = ~new_G3693gat & ~new_G3647gat;
  assign new_G3748gat = ~new_G3697gat & ~new_G3698gat;
  assign new_G3751gat = ~new_G3699gat & ~new_G1194gat;
  assign new_G3755gat = ~new_G3659gat & ~new_G3702gat;
  assign new_G3756gat = ~new_G3702gat & ~new_G1242gat;
  assign new_G3757gat = ~new_G3548gat & ~new_G3702gat;
  assign new_G3760gat = ~new_G3706gat & ~new_G567gat;
  assign new_G3764gat = ~new_G3709gat & ~new_G615gat;
  assign new_G3768gat = ~new_G3712gat & ~new_G663gat;
  assign new_G3772gat = ~new_G3715gat & ~new_G711gat;
  assign new_G3776gat = ~new_G3718gat & ~new_G759gat;
  assign new_G3780gat = ~new_G3721gat & ~new_G807gat;
  assign new_G3784gat = ~new_G3724gat & ~new_G855gat;
  assign new_G3788gat = ~new_G3727gat & ~new_G903gat;
  assign new_G3792gat = ~new_G3678gat & ~new_G3730gat;
  assign new_G3793gat = ~new_G3730gat & ~new_G951gat;
  assign new_G3794gat = ~new_G3577gat & ~new_G3730gat;
  assign new_G3797gat = ~new_G3734gat & ~new_G3735gat;
  assign new_G3800gat = ~new_G3739gat & ~new_G3736gat;
  assign new_G3804gat = ~new_G3690gat & ~new_G3742gat;
  assign new_G3805gat = ~new_G3742gat & ~new_G3687gat;
  assign new_G3806gat = ~new_G3746gat & ~new_G3747gat;
  assign new_G3809gat = ~new_G3748gat & ~new_G1146gat;
  assign new_G3813gat = ~new_G3699gat & ~new_G3751gat;
  assign new_G3814gat = ~new_G3751gat & ~new_G1194gat;
  assign new_G3815gat = ~new_G3598gat & ~new_G3751gat;
  assign new_G3818gat = ~new_G3755gat & ~new_G3756gat;
  assign new_G3821gat = ~new_G1290gat & ~new_G3757gat;
  assign new_G3825gat = ~new_G3706gat & ~new_G3760gat;
  assign new_G3826gat = ~new_G3760gat & ~new_G567gat;
  assign new_G3827gat = ~new_G3604gat & ~new_G3760gat;
  assign new_G3830gat = ~new_G3709gat & ~new_G3764gat;
  assign new_G3831gat = ~new_G3764gat & ~new_G615gat;
  assign new_G3832gat = ~new_G3608gat & ~new_G3764gat;
  assign new_G3835gat = ~new_G3712gat & ~new_G3768gat;
  assign new_G3836gat = ~new_G3768gat & ~new_G663gat;
  assign new_G3837gat = ~new_G3612gat & ~new_G3768gat;
  assign new_G3840gat = ~new_G3715gat & ~new_G3772gat;
  assign new_G3841gat = ~new_G3772gat & ~new_G711gat;
  assign new_G3842gat = ~new_G3616gat & ~new_G3772gat;
  assign new_G3845gat = ~new_G3718gat & ~new_G3776gat;
  assign new_G3846gat = ~new_G3776gat & ~new_G759gat;
  assign new_G3847gat = ~new_G3620gat & ~new_G3776gat;
  assign new_G3850gat = ~new_G3721gat & ~new_G3780gat;
  assign new_G3851gat = ~new_G3780gat & ~new_G807gat;
  assign new_G3852gat = ~new_G3624gat & ~new_G3780gat;
  assign new_G3855gat = ~new_G3724gat & ~new_G3784gat;
  assign new_G3856gat = ~new_G3784gat & ~new_G855gat;
  assign new_G3857gat = ~new_G3628gat & ~new_G3784gat;
  assign new_G3860gat = ~new_G3727gat & ~new_G3788gat;
  assign new_G3861gat = ~new_G3788gat & ~new_G903gat;
  assign new_G3862gat = ~new_G3632gat & ~new_G3788gat;
  assign new_G3865gat = ~new_G3792gat & ~new_G3793gat;
  assign new_G3868gat = ~new_G3797gat & ~new_G3794gat;
  assign new_G3872gat = ~new_G3739gat & ~new_G3800gat;
  assign new_G3873gat = ~new_G3800gat & ~new_G3736gat;
  assign new_G3874gat = ~new_G3804gat & ~new_G3805gat;
  assign new_G3877gat = ~new_G3806gat & ~new_G1098gat;
  assign new_G3881gat = ~new_G3748gat & ~new_G3809gat;
  assign new_G3882gat = ~new_G3809gat & ~new_G1146gat;
  assign new_G3883gat = ~new_G3653gat & ~new_G3809gat;
  assign new_G3886gat = ~new_G3813gat & ~new_G3814gat;
  assign new_G3889gat = ~new_G3818gat & ~new_G3815gat;
  assign new_G3893gat = ~new_G1290gat & ~new_G3821gat;
  assign new_G3894gat = ~new_G3821gat & ~new_G3757gat;
  assign G3895gat = ~new_G3825gat & ~new_G3826gat;
  assign new_G3896gat = ~new_G3830gat & ~new_G3831gat;
  assign new_G3899gat = ~new_G3835gat & ~new_G3836gat;
  assign new_G3902gat = ~new_G3840gat & ~new_G3841gat;
  assign new_G3905gat = ~new_G3845gat & ~new_G3846gat;
  assign new_G3908gat = ~new_G3850gat & ~new_G3851gat;
  assign new_G3911gat = ~new_G3855gat & ~new_G3856gat;
  assign new_G3914gat = ~new_G3860gat & ~new_G3861gat;
  assign new_G3917gat = ~new_G3865gat & ~new_G3862gat;
  assign new_G3921gat = ~new_G3797gat & ~new_G3868gat;
  assign new_G3922gat = ~new_G3868gat & ~new_G3794gat;
  assign new_G3923gat = ~new_G3872gat & ~new_G3873gat;
  assign new_G3926gat = ~new_G3874gat & ~new_G1050gat;
  assign new_G3930gat = ~new_G3806gat & ~new_G3877gat;
  assign new_G3931gat = ~new_G3877gat & ~new_G1098gat;
  assign new_G3932gat = ~new_G3693gat & ~new_G3877gat;
  assign new_G3935gat = ~new_G3881gat & ~new_G3882gat;
  assign new_G3938gat = ~new_G3886gat & ~new_G3883gat;
  assign new_G3942gat = ~new_G3818gat & ~new_G3889gat;
  assign new_G3943gat = ~new_G3889gat & ~new_G3815gat;
  assign new_G3944gat = ~new_G3893gat & ~new_G3894gat;
  assign new_G3947gat = ~new_G3896gat & ~new_G3827gat;
  assign new_G3951gat = ~new_G3899gat & ~new_G3832gat;
  assign new_G3955gat = ~new_G3902gat & ~new_G3837gat;
  assign new_G3959gat = ~new_G3905gat & ~new_G3842gat;
  assign new_G3963gat = ~new_G3908gat & ~new_G3847gat;
  assign new_G3967gat = ~new_G3911gat & ~new_G3852gat;
  assign new_G3971gat = ~new_G3914gat & ~new_G3857gat;
  assign new_G3975gat = ~new_G3865gat & ~new_G3917gat;
  assign new_G3976gat = ~new_G3917gat & ~new_G3862gat;
  assign new_G3977gat = ~new_G3921gat & ~new_G3922gat;
  assign new_G3980gat = ~new_G3923gat & ~new_G1002gat;
  assign new_G3984gat = ~new_G3874gat & ~new_G3926gat;
  assign new_G3985gat = ~new_G3926gat & ~new_G1050gat;
  assign new_G3986gat = ~new_G3742gat & ~new_G3926gat;
  assign new_G3989gat = ~new_G3930gat & ~new_G3931gat;
  assign new_G3992gat = ~new_G3935gat & ~new_G3932gat;
  assign new_G3996gat = ~new_G3886gat & ~new_G3938gat;
  assign new_G3997gat = ~new_G3938gat & ~new_G3883gat;
  assign new_G3998gat = ~new_G3942gat & ~new_G3943gat;
  assign new_G4001gat = ~new_G3944gat & ~new_G1245gat;
  assign new_G4005gat = ~new_G3896gat & ~new_G3947gat;
  assign new_G4006gat = ~new_G3947gat & ~new_G3827gat;
  assign new_G4007gat = ~new_G3899gat & ~new_G3951gat;
  assign new_G4008gat = ~new_G3951gat & ~new_G3832gat;
  assign new_G4009gat = ~new_G3902gat & ~new_G3955gat;
  assign new_G4010gat = ~new_G3955gat & ~new_G3837gat;
  assign new_G4011gat = ~new_G3905gat & ~new_G3959gat;
  assign new_G4012gat = ~new_G3959gat & ~new_G3842gat;
  assign new_G4013gat = ~new_G3908gat & ~new_G3963gat;
  assign new_G4014gat = ~new_G3963gat & ~new_G3847gat;
  assign new_G4015gat = ~new_G3911gat & ~new_G3967gat;
  assign new_G4016gat = ~new_G3967gat & ~new_G3852gat;
  assign new_G4017gat = ~new_G3914gat & ~new_G3971gat;
  assign new_G4018gat = ~new_G3971gat & ~new_G3857gat;
  assign new_G4019gat = ~new_G3975gat & ~new_G3976gat;
  assign new_G4022gat = ~new_G3977gat & ~new_G954gat;
  assign new_G4026gat = ~new_G3923gat & ~new_G3980gat;
  assign new_G4027gat = ~new_G3980gat & ~new_G1002gat;
  assign new_G4028gat = ~new_G3800gat & ~new_G3980gat;
  assign new_G4031gat = ~new_G3984gat & ~new_G3985gat;
  assign new_G4034gat = ~new_G3989gat & ~new_G3986gat;
  assign new_G4038gat = ~new_G3935gat & ~new_G3992gat;
  assign new_G4039gat = ~new_G3992gat & ~new_G3932gat;
  assign new_G4040gat = ~new_G3996gat & ~new_G3997gat;
  assign new_G4043gat = ~new_G3998gat & ~new_G1197gat;
  assign new_G4047gat = ~new_G3944gat & ~new_G4001gat;
  assign new_G4048gat = ~new_G4001gat & ~new_G1245gat;
  assign new_G4049gat = ~new_G3821gat & ~new_G4001gat;
  assign new_G4052gat = ~new_G4005gat & ~new_G4006gat;
  assign new_G4055gat = ~new_G4007gat & ~new_G4008gat;
  assign new_G4058gat = ~new_G4009gat & ~new_G4010gat;
  assign new_G4061gat = ~new_G4011gat & ~new_G4012gat;
  assign new_G4064gat = ~new_G4013gat & ~new_G4014gat;
  assign new_G4067gat = ~new_G4015gat & ~new_G4016gat;
  assign new_G4070gat = ~new_G4017gat & ~new_G4018gat;
  assign new_G4073gat = ~new_G4019gat & ~new_G906gat;
  assign new_G4077gat = ~new_G3977gat & ~new_G4022gat;
  assign new_G4078gat = ~new_G4022gat & ~new_G954gat;
  assign new_G4079gat = ~new_G3868gat & ~new_G4022gat;
  assign new_G4082gat = ~new_G4026gat & ~new_G4027gat;
  assign new_G4085gat = ~new_G4031gat & ~new_G4028gat;
  assign new_G4089gat = ~new_G3989gat & ~new_G4034gat;
  assign new_G4090gat = ~new_G4034gat & ~new_G3986gat;
  assign new_G4091gat = ~new_G4038gat & ~new_G4039gat;
  assign new_G4094gat = ~new_G4040gat & ~new_G1149gat;
  assign new_G4098gat = ~new_G3998gat & ~new_G4043gat;
  assign new_G4099gat = ~new_G4043gat & ~new_G1197gat;
  assign new_G4100gat = ~new_G3889gat & ~new_G4043gat;
  assign new_G4103gat = ~new_G4047gat & ~new_G4048gat;
  assign new_G4106gat = ~new_G1293gat & ~new_G4049gat;
  assign new_G4110gat = ~new_G4052gat & ~new_G570gat;
  assign new_G4114gat = ~new_G4055gat & ~new_G618gat;
  assign new_G4118gat = ~new_G4058gat & ~new_G666gat;
  assign new_G4122gat = ~new_G4061gat & ~new_G714gat;
  assign new_G4126gat = ~new_G4064gat & ~new_G762gat;
  assign new_G4130gat = ~new_G4067gat & ~new_G810gat;
  assign new_G4134gat = ~new_G4070gat & ~new_G858gat;
  assign new_G4138gat = ~new_G4019gat & ~new_G4073gat;
  assign new_G4139gat = ~new_G4073gat & ~new_G906gat;
  assign new_G4140gat = ~new_G3917gat & ~new_G4073gat;
  assign new_G4143gat = ~new_G4077gat & ~new_G4078gat;
  assign new_G4146gat = ~new_G4082gat & ~new_G4079gat;
  assign new_G4150gat = ~new_G4031gat & ~new_G4085gat;
  assign new_G4151gat = ~new_G4085gat & ~new_G4028gat;
  assign new_G4152gat = ~new_G4089gat & ~new_G4090gat;
  assign new_G4155gat = ~new_G4091gat & ~new_G1101gat;
  assign new_G4159gat = ~new_G4040gat & ~new_G4094gat;
  assign new_G4160gat = ~new_G4094gat & ~new_G1149gat;
  assign new_G4161gat = ~new_G3938gat & ~new_G4094gat;
  assign new_G4164gat = ~new_G4098gat & ~new_G4099gat;
  assign new_G4167gat = ~new_G4103gat & ~new_G4100gat;
  assign new_G4171gat = ~new_G1293gat & ~new_G4106gat;
  assign new_G4172gat = ~new_G4106gat & ~new_G4049gat;
  assign new_G4173gat = ~new_G4052gat & ~new_G4110gat;
  assign new_G4174gat = ~new_G4110gat & ~new_G570gat;
  assign new_G4175gat = ~new_G3947gat & ~new_G4110gat;
  assign new_G4178gat = ~new_G4055gat & ~new_G4114gat;
  assign new_G4179gat = ~new_G4114gat & ~new_G618gat;
  assign new_G4180gat = ~new_G3951gat & ~new_G4114gat;
  assign new_G4183gat = ~new_G4058gat & ~new_G4118gat;
  assign new_G4184gat = ~new_G4118gat & ~new_G666gat;
  assign new_G4185gat = ~new_G3955gat & ~new_G4118gat;
  assign new_G4188gat = ~new_G4061gat & ~new_G4122gat;
  assign new_G4189gat = ~new_G4122gat & ~new_G714gat;
  assign new_G4190gat = ~new_G3959gat & ~new_G4122gat;
  assign new_G4193gat = ~new_G4064gat & ~new_G4126gat;
  assign new_G4194gat = ~new_G4126gat & ~new_G762gat;
  assign new_G4195gat = ~new_G3963gat & ~new_G4126gat;
  assign new_G4198gat = ~new_G4067gat & ~new_G4130gat;
  assign new_G4199gat = ~new_G4130gat & ~new_G810gat;
  assign new_G4200gat = ~new_G3967gat & ~new_G4130gat;
  assign new_G4203gat = ~new_G4070gat & ~new_G4134gat;
  assign new_G4204gat = ~new_G4134gat & ~new_G858gat;
  assign new_G4205gat = ~new_G3971gat & ~new_G4134gat;
  assign new_G4208gat = ~new_G4138gat & ~new_G4139gat;
  assign new_G4211gat = ~new_G4143gat & ~new_G4140gat;
  assign new_G4215gat = ~new_G4082gat & ~new_G4146gat;
  assign new_G4216gat = ~new_G4146gat & ~new_G4079gat;
  assign new_G4217gat = ~new_G4150gat & ~new_G4151gat;
  assign new_G4220gat = ~new_G4152gat & ~new_G1053gat;
  assign new_G4224gat = ~new_G4091gat & ~new_G4155gat;
  assign new_G4225gat = ~new_G4155gat & ~new_G1101gat;
  assign new_G4226gat = ~new_G3992gat & ~new_G4155gat;
  assign new_G4229gat = ~new_G4159gat & ~new_G4160gat;
  assign new_G4232gat = ~new_G4164gat & ~new_G4161gat;
  assign new_G4236gat = ~new_G4103gat & ~new_G4167gat;
  assign new_G4237gat = ~new_G4167gat & ~new_G4100gat;
  assign new_G4238gat = ~new_G4171gat & ~new_G4172gat;
  assign G4241gat = ~new_G4173gat & ~new_G4174gat;
  assign new_G4242gat = ~new_G4178gat & ~new_G4179gat;
  assign new_G4245gat = ~new_G4183gat & ~new_G4184gat;
  assign new_G4248gat = ~new_G4188gat & ~new_G4189gat;
  assign new_G4251gat = ~new_G4193gat & ~new_G4194gat;
  assign new_G4254gat = ~new_G4198gat & ~new_G4199gat;
  assign new_G4257gat = ~new_G4203gat & ~new_G4204gat;
  assign new_G4260gat = ~new_G4208gat & ~new_G4205gat;
  assign new_G4264gat = ~new_G4143gat & ~new_G4211gat;
  assign new_G4265gat = ~new_G4211gat & ~new_G4140gat;
  assign new_G4266gat = ~new_G4215gat & ~new_G4216gat;
  assign new_G4269gat = ~new_G4217gat & ~new_G1005gat;
  assign new_G4273gat = ~new_G4152gat & ~new_G4220gat;
  assign new_G4274gat = ~new_G4220gat & ~new_G1053gat;
  assign new_G4275gat = ~new_G4034gat & ~new_G4220gat;
  assign new_G4278gat = ~new_G4224gat & ~new_G4225gat;
  assign new_G4281gat = ~new_G4229gat & ~new_G4226gat;
  assign new_G4285gat = ~new_G4164gat & ~new_G4232gat;
  assign new_G4286gat = ~new_G4232gat & ~new_G4161gat;
  assign new_G4287gat = ~new_G4236gat & ~new_G4237gat;
  assign new_G4290gat = ~new_G4238gat & ~new_G1248gat;
  assign new_G4294gat = ~new_G4242gat & ~new_G4175gat;
  assign new_G4298gat = ~new_G4245gat & ~new_G4180gat;
  assign new_G4302gat = ~new_G4248gat & ~new_G4185gat;
  assign new_G4306gat = ~new_G4251gat & ~new_G4190gat;
  assign new_G4310gat = ~new_G4254gat & ~new_G4195gat;
  assign new_G4314gat = ~new_G4257gat & ~new_G4200gat;
  assign new_G4318gat = ~new_G4208gat & ~new_G4260gat;
  assign new_G4319gat = ~new_G4260gat & ~new_G4205gat;
  assign new_G4320gat = ~new_G4264gat & ~new_G4265gat;
  assign new_G4323gat = ~new_G4266gat & ~new_G957gat;
  assign new_G4327gat = ~new_G4217gat & ~new_G4269gat;
  assign new_G4328gat = ~new_G4269gat & ~new_G1005gat;
  assign new_G4329gat = ~new_G4085gat & ~new_G4269gat;
  assign new_G4332gat = ~new_G4273gat & ~new_G4274gat;
  assign new_G4335gat = ~new_G4278gat & ~new_G4275gat;
  assign new_G4339gat = ~new_G4229gat & ~new_G4281gat;
  assign new_G4340gat = ~new_G4281gat & ~new_G4226gat;
  assign new_G4341gat = ~new_G4285gat & ~new_G4286gat;
  assign new_G4344gat = ~new_G4287gat & ~new_G1200gat;
  assign new_G4348gat = ~new_G4238gat & ~new_G4290gat;
  assign new_G4349gat = ~new_G4290gat & ~new_G1248gat;
  assign new_G4350gat = ~new_G4106gat & ~new_G4290gat;
  assign new_G4353gat = ~new_G4242gat & ~new_G4294gat;
  assign new_G4354gat = ~new_G4294gat & ~new_G4175gat;
  assign new_G4355gat = ~new_G4245gat & ~new_G4298gat;
  assign new_G4356gat = ~new_G4298gat & ~new_G4180gat;
  assign new_G4357gat = ~new_G4248gat & ~new_G4302gat;
  assign new_G4358gat = ~new_G4302gat & ~new_G4185gat;
  assign new_G4359gat = ~new_G4251gat & ~new_G4306gat;
  assign new_G4360gat = ~new_G4306gat & ~new_G4190gat;
  assign new_G4361gat = ~new_G4254gat & ~new_G4310gat;
  assign new_G4362gat = ~new_G4310gat & ~new_G4195gat;
  assign new_G4363gat = ~new_G4257gat & ~new_G4314gat;
  assign new_G4364gat = ~new_G4314gat & ~new_G4200gat;
  assign new_G4365gat = ~new_G4318gat & ~new_G4319gat;
  assign new_G4368gat = ~new_G4320gat & ~new_G909gat;
  assign new_G4372gat = ~new_G4266gat & ~new_G4323gat;
  assign new_G4373gat = ~new_G4323gat & ~new_G957gat;
  assign new_G4374gat = ~new_G4146gat & ~new_G4323gat;
  assign new_G4377gat = ~new_G4327gat & ~new_G4328gat;
  assign new_G4380gat = ~new_G4332gat & ~new_G4329gat;
  assign new_G4384gat = ~new_G4278gat & ~new_G4335gat;
  assign new_G4385gat = ~new_G4335gat & ~new_G4275gat;
  assign new_G4386gat = ~new_G4339gat & ~new_G4340gat;
  assign new_G4389gat = ~new_G4341gat & ~new_G1152gat;
  assign new_G4393gat = ~new_G4287gat & ~new_G4344gat;
  assign new_G4394gat = ~new_G4344gat & ~new_G1200gat;
  assign new_G4395gat = ~new_G4167gat & ~new_G4344gat;
  assign new_G4398gat = ~new_G4348gat & ~new_G4349gat;
  assign new_G4401gat = ~new_G1296gat & ~new_G4350gat;
  assign new_G4405gat = ~new_G4353gat & ~new_G4354gat;
  assign new_G4408gat = ~new_G4355gat & ~new_G4356gat;
  assign new_G4411gat = ~new_G4357gat & ~new_G4358gat;
  assign new_G4414gat = ~new_G4359gat & ~new_G4360gat;
  assign new_G4417gat = ~new_G4361gat & ~new_G4362gat;
  assign new_G4420gat = ~new_G4363gat & ~new_G4364gat;
  assign new_G4423gat = ~new_G4365gat & ~new_G861gat;
  assign new_G4427gat = ~new_G4320gat & ~new_G4368gat;
  assign new_G4428gat = ~new_G4368gat & ~new_G909gat;
  assign new_G4429gat = ~new_G4211gat & ~new_G4368gat;
  assign new_G4432gat = ~new_G4372gat & ~new_G4373gat;
  assign new_G4435gat = ~new_G4377gat & ~new_G4374gat;
  assign new_G4439gat = ~new_G4332gat & ~new_G4380gat;
  assign new_G4440gat = ~new_G4380gat & ~new_G4329gat;
  assign new_G4441gat = ~new_G4384gat & ~new_G4385gat;
  assign new_G4444gat = ~new_G4386gat & ~new_G1104gat;
  assign new_G4448gat = ~new_G4341gat & ~new_G4389gat;
  assign new_G4449gat = ~new_G4389gat & ~new_G1152gat;
  assign new_G4450gat = ~new_G4232gat & ~new_G4389gat;
  assign new_G4453gat = ~new_G4393gat & ~new_G4394gat;
  assign new_G4456gat = ~new_G4398gat & ~new_G4395gat;
  assign new_G4460gat = ~new_G1296gat & ~new_G4401gat;
  assign new_G4461gat = ~new_G4401gat & ~new_G4350gat;
  assign new_G4462gat = ~new_G4405gat & ~new_G573gat;
  assign new_G4466gat = ~new_G4408gat & ~new_G621gat;
  assign new_G4470gat = ~new_G4411gat & ~new_G669gat;
  assign new_G4474gat = ~new_G4414gat & ~new_G717gat;
  assign new_G4478gat = ~new_G4417gat & ~new_G765gat;
  assign new_G4482gat = ~new_G4420gat & ~new_G813gat;
  assign new_G4486gat = ~new_G4365gat & ~new_G4423gat;
  assign new_G4487gat = ~new_G4423gat & ~new_G861gat;
  assign new_G4488gat = ~new_G4260gat & ~new_G4423gat;
  assign new_G4491gat = ~new_G4427gat & ~new_G4428gat;
  assign new_G4494gat = ~new_G4432gat & ~new_G4429gat;
  assign new_G4498gat = ~new_G4377gat & ~new_G4435gat;
  assign new_G4499gat = ~new_G4435gat & ~new_G4374gat;
  assign new_G4500gat = ~new_G4439gat & ~new_G4440gat;
  assign new_G4503gat = ~new_G4441gat & ~new_G1056gat;
  assign new_G4507gat = ~new_G4386gat & ~new_G4444gat;
  assign new_G4508gat = ~new_G4444gat & ~new_G1104gat;
  assign new_G4509gat = ~new_G4281gat & ~new_G4444gat;
  assign new_G4512gat = ~new_G4448gat & ~new_G4449gat;
  assign new_G4515gat = ~new_G4453gat & ~new_G4450gat;
  assign new_G4519gat = ~new_G4398gat & ~new_G4456gat;
  assign new_G4520gat = ~new_G4456gat & ~new_G4395gat;
  assign new_G4521gat = ~new_G4460gat & ~new_G4461gat;
  assign new_G4524gat = ~new_G4405gat & ~new_G4462gat;
  assign new_G4525gat = ~new_G4462gat & ~new_G573gat;
  assign new_G4526gat = ~new_G4294gat & ~new_G4462gat;
  assign new_G4529gat = ~new_G4408gat & ~new_G4466gat;
  assign new_G4530gat = ~new_G4466gat & ~new_G621gat;
  assign new_G4531gat = ~new_G4298gat & ~new_G4466gat;
  assign new_G4534gat = ~new_G4411gat & ~new_G4470gat;
  assign new_G4535gat = ~new_G4470gat & ~new_G669gat;
  assign new_G4536gat = ~new_G4302gat & ~new_G4470gat;
  assign new_G4539gat = ~new_G4414gat & ~new_G4474gat;
  assign new_G4540gat = ~new_G4474gat & ~new_G717gat;
  assign new_G4541gat = ~new_G4306gat & ~new_G4474gat;
  assign new_G4544gat = ~new_G4417gat & ~new_G4478gat;
  assign new_G4545gat = ~new_G4478gat & ~new_G765gat;
  assign new_G4546gat = ~new_G4310gat & ~new_G4478gat;
  assign new_G4549gat = ~new_G4420gat & ~new_G4482gat;
  assign new_G4550gat = ~new_G4482gat & ~new_G813gat;
  assign new_G4551gat = ~new_G4314gat & ~new_G4482gat;
  assign new_G4554gat = ~new_G4486gat & ~new_G4487gat;
  assign new_G4557gat = ~new_G4491gat & ~new_G4488gat;
  assign new_G4561gat = ~new_G4432gat & ~new_G4494gat;
  assign new_G4562gat = ~new_G4494gat & ~new_G4429gat;
  assign new_G4563gat = ~new_G4498gat & ~new_G4499gat;
  assign new_G4566gat = ~new_G4500gat & ~new_G1008gat;
  assign new_G4570gat = ~new_G4441gat & ~new_G4503gat;
  assign new_G4571gat = ~new_G4503gat & ~new_G1056gat;
  assign new_G4572gat = ~new_G4335gat & ~new_G4503gat;
  assign new_G4575gat = ~new_G4507gat & ~new_G4508gat;
  assign new_G4578gat = ~new_G4512gat & ~new_G4509gat;
  assign new_G4582gat = ~new_G4453gat & ~new_G4515gat;
  assign new_G4583gat = ~new_G4515gat & ~new_G4450gat;
  assign new_G4584gat = ~new_G4519gat & ~new_G4520gat;
  assign new_G4587gat = ~new_G4521gat & ~new_G1251gat;
  assign G4591gat = ~new_G4524gat & ~new_G4525gat;
  assign new_G4592gat = ~new_G4529gat & ~new_G4530gat;
  assign new_G4595gat = ~new_G4534gat & ~new_G4535gat;
  assign new_G4598gat = ~new_G4539gat & ~new_G4540gat;
  assign new_G4601gat = ~new_G4544gat & ~new_G4545gat;
  assign new_G4604gat = ~new_G4549gat & ~new_G4550gat;
  assign new_G4607gat = ~new_G4554gat & ~new_G4551gat;
  assign new_G4611gat = ~new_G4491gat & ~new_G4557gat;
  assign new_G4612gat = ~new_G4557gat & ~new_G4488gat;
  assign new_G4613gat = ~new_G4561gat & ~new_G4562gat;
  assign new_G4616gat = ~new_G4563gat & ~new_G960gat;
  assign new_G4620gat = ~new_G4500gat & ~new_G4566gat;
  assign new_G4621gat = ~new_G4566gat & ~new_G1008gat;
  assign new_G4622gat = ~new_G4380gat & ~new_G4566gat;
  assign new_G4625gat = ~new_G4570gat & ~new_G4571gat;
  assign new_G4628gat = ~new_G4575gat & ~new_G4572gat;
  assign new_G4632gat = ~new_G4512gat & ~new_G4578gat;
  assign new_G4633gat = ~new_G4578gat & ~new_G4509gat;
  assign new_G4634gat = ~new_G4582gat & ~new_G4583gat;
  assign new_G4637gat = ~new_G4584gat & ~new_G1203gat;
  assign new_G4641gat = ~new_G4521gat & ~new_G4587gat;
  assign new_G4642gat = ~new_G4587gat & ~new_G1251gat;
  assign new_G4643gat = ~new_G4401gat & ~new_G4587gat;
  assign new_G4646gat = ~new_G4592gat & ~new_G4526gat;
  assign new_G4650gat = ~new_G4595gat & ~new_G4531gat;
  assign new_G4654gat = ~new_G4598gat & ~new_G4536gat;
  assign new_G4658gat = ~new_G4601gat & ~new_G4541gat;
  assign new_G4662gat = ~new_G4604gat & ~new_G4546gat;
  assign new_G4666gat = ~new_G4554gat & ~new_G4607gat;
  assign new_G4667gat = ~new_G4607gat & ~new_G4551gat;
  assign new_G4668gat = ~new_G4611gat & ~new_G4612gat;
  assign new_G4671gat = ~new_G4613gat & ~new_G912gat;
  assign new_G4675gat = ~new_G4563gat & ~new_G4616gat;
  assign new_G4676gat = ~new_G4616gat & ~new_G960gat;
  assign new_G4677gat = ~new_G4435gat & ~new_G4616gat;
  assign new_G4680gat = ~new_G4620gat & ~new_G4621gat;
  assign new_G4683gat = ~new_G4625gat & ~new_G4622gat;
  assign new_G4687gat = ~new_G4575gat & ~new_G4628gat;
  assign new_G4688gat = ~new_G4628gat & ~new_G4572gat;
  assign new_G4689gat = ~new_G4632gat & ~new_G4633gat;
  assign new_G4692gat = ~new_G4634gat & ~new_G1155gat;
  assign new_G4696gat = ~new_G4584gat & ~new_G4637gat;
  assign new_G4697gat = ~new_G4637gat & ~new_G1203gat;
  assign new_G4698gat = ~new_G4456gat & ~new_G4637gat;
  assign new_G4701gat = ~new_G4641gat & ~new_G4642gat;
  assign new_G4704gat = ~new_G1299gat & ~new_G4643gat;
  assign new_G4708gat = ~new_G4592gat & ~new_G4646gat;
  assign new_G4709gat = ~new_G4646gat & ~new_G4526gat;
  assign new_G4710gat = ~new_G4595gat & ~new_G4650gat;
  assign new_G4711gat = ~new_G4650gat & ~new_G4531gat;
  assign new_G4712gat = ~new_G4598gat & ~new_G4654gat;
  assign new_G4713gat = ~new_G4654gat & ~new_G4536gat;
  assign new_G4714gat = ~new_G4601gat & ~new_G4658gat;
  assign new_G4715gat = ~new_G4658gat & ~new_G4541gat;
  assign new_G4716gat = ~new_G4604gat & ~new_G4662gat;
  assign new_G4717gat = ~new_G4662gat & ~new_G4546gat;
  assign new_G4718gat = ~new_G4666gat & ~new_G4667gat;
  assign new_G4721gat = ~new_G4668gat & ~new_G864gat;
  assign new_G4725gat = ~new_G4613gat & ~new_G4671gat;
  assign new_G4726gat = ~new_G4671gat & ~new_G912gat;
  assign new_G4727gat = ~new_G4494gat & ~new_G4671gat;
  assign new_G4730gat = ~new_G4675gat & ~new_G4676gat;
  assign new_G4733gat = ~new_G4680gat & ~new_G4677gat;
  assign new_G4737gat = ~new_G4625gat & ~new_G4683gat;
  assign new_G4738gat = ~new_G4683gat & ~new_G4622gat;
  assign new_G4739gat = ~new_G4687gat & ~new_G4688gat;
  assign new_G4742gat = ~new_G4689gat & ~new_G1107gat;
  assign new_G4746gat = ~new_G4634gat & ~new_G4692gat;
  assign new_G4747gat = ~new_G4692gat & ~new_G1155gat;
  assign new_G4748gat = ~new_G4515gat & ~new_G4692gat;
  assign new_G4751gat = ~new_G4696gat & ~new_G4697gat;
  assign new_G4754gat = ~new_G4701gat & ~new_G4698gat;
  assign new_G4758gat = ~new_G1299gat & ~new_G4704gat;
  assign new_G4759gat = ~new_G4704gat & ~new_G4643gat;
  assign new_G4760gat = ~new_G4708gat & ~new_G4709gat;
  assign new_G4763gat = ~new_G4710gat & ~new_G4711gat;
  assign new_G4766gat = ~new_G4712gat & ~new_G4713gat;
  assign new_G4769gat = ~new_G4714gat & ~new_G4715gat;
  assign new_G4772gat = ~new_G4716gat & ~new_G4717gat;
  assign new_G4775gat = ~new_G4718gat & ~new_G816gat;
  assign new_G4779gat = ~new_G4668gat & ~new_G4721gat;
  assign new_G4780gat = ~new_G4721gat & ~new_G864gat;
  assign new_G4781gat = ~new_G4557gat & ~new_G4721gat;
  assign new_G4784gat = ~new_G4725gat & ~new_G4726gat;
  assign new_G4787gat = ~new_G4730gat & ~new_G4727gat;
  assign new_G4791gat = ~new_G4680gat & ~new_G4733gat;
  assign new_G4792gat = ~new_G4733gat & ~new_G4677gat;
  assign new_G4793gat = ~new_G4737gat & ~new_G4738gat;
  assign new_G4796gat = ~new_G4739gat & ~new_G1059gat;
  assign new_G4800gat = ~new_G4689gat & ~new_G4742gat;
  assign new_G4801gat = ~new_G4742gat & ~new_G1107gat;
  assign new_G4802gat = ~new_G4578gat & ~new_G4742gat;
  assign new_G4805gat = ~new_G4746gat & ~new_G4747gat;
  assign new_G4808gat = ~new_G4751gat & ~new_G4748gat;
  assign new_G4812gat = ~new_G4701gat & ~new_G4754gat;
  assign new_G4813gat = ~new_G4754gat & ~new_G4698gat;
  assign new_G4814gat = ~new_G4758gat & ~new_G4759gat;
  assign new_G4817gat = ~new_G4760gat & ~new_G576gat;
  assign new_G4821gat = ~new_G4763gat & ~new_G624gat;
  assign new_G4825gat = ~new_G4766gat & ~new_G672gat;
  assign new_G4829gat = ~new_G4769gat & ~new_G720gat;
  assign new_G4833gat = ~new_G4772gat & ~new_G768gat;
  assign new_G4837gat = ~new_G4718gat & ~new_G4775gat;
  assign new_G4838gat = ~new_G4775gat & ~new_G816gat;
  assign new_G4839gat = ~new_G4607gat & ~new_G4775gat;
  assign new_G4842gat = ~new_G4779gat & ~new_G4780gat;
  assign new_G4845gat = ~new_G4784gat & ~new_G4781gat;
  assign new_G4849gat = ~new_G4730gat & ~new_G4787gat;
  assign new_G4850gat = ~new_G4787gat & ~new_G4727gat;
  assign new_G4851gat = ~new_G4791gat & ~new_G4792gat;
  assign new_G4854gat = ~new_G4793gat & ~new_G1011gat;
  assign new_G4858gat = ~new_G4739gat & ~new_G4796gat;
  assign new_G4859gat = ~new_G4796gat & ~new_G1059gat;
  assign new_G4860gat = ~new_G4628gat & ~new_G4796gat;
  assign new_G4863gat = ~new_G4800gat & ~new_G4801gat;
  assign new_G4866gat = ~new_G4805gat & ~new_G4802gat;
  assign new_G4870gat = ~new_G4751gat & ~new_G4808gat;
  assign new_G4871gat = ~new_G4808gat & ~new_G4748gat;
  assign new_G4872gat = ~new_G4812gat & ~new_G4813gat;
  assign new_G4875gat = ~new_G4814gat & ~new_G1254gat;
  assign new_G4879gat = ~new_G4760gat & ~new_G4817gat;
  assign new_G4880gat = ~new_G4817gat & ~new_G576gat;
  assign new_G4881gat = ~new_G4646gat & ~new_G4817gat;
  assign new_G4884gat = ~new_G4763gat & ~new_G4821gat;
  assign new_G4885gat = ~new_G4821gat & ~new_G624gat;
  assign new_G4886gat = ~new_G4650gat & ~new_G4821gat;
  assign new_G4889gat = ~new_G4766gat & ~new_G4825gat;
  assign new_G4890gat = ~new_G4825gat & ~new_G672gat;
  assign new_G4891gat = ~new_G4654gat & ~new_G4825gat;
  assign new_G4894gat = ~new_G4769gat & ~new_G4829gat;
  assign new_G4895gat = ~new_G4829gat & ~new_G720gat;
  assign new_G4896gat = ~new_G4658gat & ~new_G4829gat;
  assign new_G4899gat = ~new_G4772gat & ~new_G4833gat;
  assign new_G4900gat = ~new_G4833gat & ~new_G768gat;
  assign new_G4901gat = ~new_G4662gat & ~new_G4833gat;
  assign new_G4904gat = ~new_G4837gat & ~new_G4838gat;
  assign new_G4907gat = ~new_G4842gat & ~new_G4839gat;
  assign new_G4911gat = ~new_G4784gat & ~new_G4845gat;
  assign new_G4912gat = ~new_G4845gat & ~new_G4781gat;
  assign new_G4913gat = ~new_G4849gat & ~new_G4850gat;
  assign new_G4916gat = ~new_G4851gat & ~new_G963gat;
  assign new_G4920gat = ~new_G4793gat & ~new_G4854gat;
  assign new_G4921gat = ~new_G4854gat & ~new_G1011gat;
  assign new_G4922gat = ~new_G4683gat & ~new_G4854gat;
  assign new_G4925gat = ~new_G4858gat & ~new_G4859gat;
  assign new_G4928gat = ~new_G4863gat & ~new_G4860gat;
  assign new_G4932gat = ~new_G4805gat & ~new_G4866gat;
  assign new_G4933gat = ~new_G4866gat & ~new_G4802gat;
  assign new_G4934gat = ~new_G4870gat & ~new_G4871gat;
  assign new_G4937gat = ~new_G4872gat & ~new_G1206gat;
  assign new_G4941gat = ~new_G4814gat & ~new_G4875gat;
  assign new_G4942gat = ~new_G4875gat & ~new_G1254gat;
  assign new_G4943gat = ~new_G4704gat & ~new_G4875gat;
  assign G4946gat = ~new_G4879gat & ~new_G4880gat;
  assign new_G4947gat = ~new_G4884gat & ~new_G4885gat;
  assign new_G4950gat = ~new_G4889gat & ~new_G4890gat;
  assign new_G4953gat = ~new_G4894gat & ~new_G4895gat;
  assign new_G4956gat = ~new_G4899gat & ~new_G4900gat;
  assign new_G4959gat = ~new_G4904gat & ~new_G4901gat;
  assign new_G4963gat = ~new_G4842gat & ~new_G4907gat;
  assign new_G4964gat = ~new_G4907gat & ~new_G4839gat;
  assign new_G4965gat = ~new_G4911gat & ~new_G4912gat;
  assign new_G4968gat = ~new_G4913gat & ~new_G915gat;
  assign new_G4972gat = ~new_G4851gat & ~new_G4916gat;
  assign new_G4973gat = ~new_G4916gat & ~new_G963gat;
  assign new_G4974gat = ~new_G4733gat & ~new_G4916gat;
  assign new_G4977gat = ~new_G4920gat & ~new_G4921gat;
  assign new_G4980gat = ~new_G4925gat & ~new_G4922gat;
  assign new_G4984gat = ~new_G4863gat & ~new_G4928gat;
  assign new_G4985gat = ~new_G4928gat & ~new_G4860gat;
  assign new_G4986gat = ~new_G4932gat & ~new_G4933gat;
  assign new_G4989gat = ~new_G4934gat & ~new_G1158gat;
  assign new_G4993gat = ~new_G4872gat & ~new_G4937gat;
  assign new_G4994gat = ~new_G4937gat & ~new_G1206gat;
  assign new_G4995gat = ~new_G4754gat & ~new_G4937gat;
  assign new_G4998gat = ~new_G4941gat & ~new_G4942gat;
  assign new_G5001gat = ~new_G1302gat & ~new_G4943gat;
  assign new_G5005gat = ~new_G4947gat & ~new_G4881gat;
  assign new_G5009gat = ~new_G4950gat & ~new_G4886gat;
  assign new_G5013gat = ~new_G4953gat & ~new_G4891gat;
  assign new_G5017gat = ~new_G4956gat & ~new_G4896gat;
  assign new_G5021gat = ~new_G4904gat & ~new_G4959gat;
  assign new_G5022gat = ~new_G4959gat & ~new_G4901gat;
  assign new_G5023gat = ~new_G4963gat & ~new_G4964gat;
  assign new_G5026gat = ~new_G4965gat & ~new_G867gat;
  assign new_G5030gat = ~new_G4913gat & ~new_G4968gat;
  assign new_G5031gat = ~new_G4968gat & ~new_G915gat;
  assign new_G5032gat = ~new_G4787gat & ~new_G4968gat;
  assign new_G5035gat = ~new_G4972gat & ~new_G4973gat;
  assign new_G5038gat = ~new_G4977gat & ~new_G4974gat;
  assign new_G5042gat = ~new_G4925gat & ~new_G4980gat;
  assign new_G5043gat = ~new_G4980gat & ~new_G4922gat;
  assign new_G5044gat = ~new_G4984gat & ~new_G4985gat;
  assign new_G5047gat = ~new_G4986gat & ~new_G1110gat;
  assign new_G5051gat = ~new_G4934gat & ~new_G4989gat;
  assign new_G5052gat = ~new_G4989gat & ~new_G1158gat;
  assign new_G5053gat = ~new_G4808gat & ~new_G4989gat;
  assign new_G5056gat = ~new_G4993gat & ~new_G4994gat;
  assign new_G5059gat = ~new_G4998gat & ~new_G4995gat;
  assign new_G5063gat = ~new_G1302gat & ~new_G5001gat;
  assign new_G5064gat = ~new_G5001gat & ~new_G4943gat;
  assign new_G5065gat = ~new_G4947gat & ~new_G5005gat;
  assign new_G5066gat = ~new_G5005gat & ~new_G4881gat;
  assign new_G5067gat = ~new_G4950gat & ~new_G5009gat;
  assign new_G5068gat = ~new_G5009gat & ~new_G4886gat;
  assign new_G5069gat = ~new_G4953gat & ~new_G5013gat;
  assign new_G5070gat = ~new_G5013gat & ~new_G4891gat;
  assign new_G5071gat = ~new_G4956gat & ~new_G5017gat;
  assign new_G5072gat = ~new_G5017gat & ~new_G4896gat;
  assign new_G5073gat = ~new_G5021gat & ~new_G5022gat;
  assign new_G5076gat = ~new_G5023gat & ~new_G819gat;
  assign new_G5080gat = ~new_G4965gat & ~new_G5026gat;
  assign new_G5081gat = ~new_G5026gat & ~new_G867gat;
  assign new_G5082gat = ~new_G4845gat & ~new_G5026gat;
  assign new_G5085gat = ~new_G5030gat & ~new_G5031gat;
  assign new_G5088gat = ~new_G5035gat & ~new_G5032gat;
  assign new_G5092gat = ~new_G4977gat & ~new_G5038gat;
  assign new_G5093gat = ~new_G5038gat & ~new_G4974gat;
  assign new_G5094gat = ~new_G5042gat & ~new_G5043gat;
  assign new_G5097gat = ~new_G5044gat & ~new_G1062gat;
  assign new_G5101gat = ~new_G4986gat & ~new_G5047gat;
  assign new_G5102gat = ~new_G5047gat & ~new_G1110gat;
  assign new_G5103gat = ~new_G4866gat & ~new_G5047gat;
  assign new_G5106gat = ~new_G5051gat & ~new_G5052gat;
  assign new_G5109gat = ~new_G5056gat & ~new_G5053gat;
  assign new_G5113gat = ~new_G4998gat & ~new_G5059gat;
  assign new_G5114gat = ~new_G5059gat & ~new_G4995gat;
  assign new_G5115gat = ~new_G5063gat & ~new_G5064gat;
  assign new_G5118gat = ~new_G5065gat & ~new_G5066gat;
  assign new_G5121gat = ~new_G5067gat & ~new_G5068gat;
  assign new_G5124gat = ~new_G5069gat & ~new_G5070gat;
  assign new_G5127gat = ~new_G5071gat & ~new_G5072gat;
  assign new_G5130gat = ~new_G5073gat & ~new_G771gat;
  assign new_G5134gat = ~new_G5023gat & ~new_G5076gat;
  assign new_G5135gat = ~new_G5076gat & ~new_G819gat;
  assign new_G5136gat = ~new_G4907gat & ~new_G5076gat;
  assign new_G5139gat = ~new_G5080gat & ~new_G5081gat;
  assign new_G5142gat = ~new_G5085gat & ~new_G5082gat;
  assign new_G5146gat = ~new_G5035gat & ~new_G5088gat;
  assign new_G5147gat = ~new_G5088gat & ~new_G5032gat;
  assign new_G5148gat = ~new_G5092gat & ~new_G5093gat;
  assign new_G5151gat = ~new_G5094gat & ~new_G1014gat;
  assign new_G5155gat = ~new_G5044gat & ~new_G5097gat;
  assign new_G5156gat = ~new_G5097gat & ~new_G1062gat;
  assign new_G5157gat = ~new_G4928gat & ~new_G5097gat;
  assign new_G5160gat = ~new_G5101gat & ~new_G5102gat;
  assign new_G5163gat = ~new_G5106gat & ~new_G5103gat;
  assign new_G5167gat = ~new_G5056gat & ~new_G5109gat;
  assign new_G5168gat = ~new_G5109gat & ~new_G5053gat;
  assign new_G5169gat = ~new_G5113gat & ~new_G5114gat;
  assign new_G5172gat = ~new_G5115gat & ~new_G1257gat;
  assign new_G5176gat = ~new_G5118gat & ~new_G579gat;
  assign new_G5180gat = ~new_G5121gat & ~new_G627gat;
  assign new_G5184gat = ~new_G5124gat & ~new_G675gat;
  assign new_G5188gat = ~new_G5127gat & ~new_G723gat;
  assign new_G5192gat = ~new_G5073gat & ~new_G5130gat;
  assign new_G5193gat = ~new_G5130gat & ~new_G771gat;
  assign new_G5194gat = ~new_G4959gat & ~new_G5130gat;
  assign new_G5197gat = ~new_G5134gat & ~new_G5135gat;
  assign new_G5200gat = ~new_G5139gat & ~new_G5136gat;
  assign new_G5204gat = ~new_G5085gat & ~new_G5142gat;
  assign new_G5205gat = ~new_G5142gat & ~new_G5082gat;
  assign new_G5206gat = ~new_G5146gat & ~new_G5147gat;
  assign new_G5209gat = ~new_G5148gat & ~new_G966gat;
  assign new_G5213gat = ~new_G5094gat & ~new_G5151gat;
  assign new_G5214gat = ~new_G5151gat & ~new_G1014gat;
  assign new_G5215gat = ~new_G4980gat & ~new_G5151gat;
  assign new_G5218gat = ~new_G5155gat & ~new_G5156gat;
  assign new_G5221gat = ~new_G5160gat & ~new_G5157gat;
  assign new_G5225gat = ~new_G5106gat & ~new_G5163gat;
  assign new_G5226gat = ~new_G5163gat & ~new_G5103gat;
  assign new_G5227gat = ~new_G5167gat & ~new_G5168gat;
  assign new_G5230gat = ~new_G5169gat & ~new_G1209gat;
  assign new_G5234gat = ~new_G5115gat & ~new_G5172gat;
  assign new_G5235gat = ~new_G5172gat & ~new_G1257gat;
  assign new_G5236gat = ~new_G5001gat & ~new_G5172gat;
  assign new_G5239gat = ~new_G5118gat & ~new_G5176gat;
  assign new_G5240gat = ~new_G5176gat & ~new_G579gat;
  assign new_G5241gat = ~new_G5005gat & ~new_G5176gat;
  assign new_G5244gat = ~new_G5121gat & ~new_G5180gat;
  assign new_G5245gat = ~new_G5180gat & ~new_G627gat;
  assign new_G5246gat = ~new_G5009gat & ~new_G5180gat;
  assign new_G5249gat = ~new_G5124gat & ~new_G5184gat;
  assign new_G5250gat = ~new_G5184gat & ~new_G675gat;
  assign new_G5251gat = ~new_G5013gat & ~new_G5184gat;
  assign new_G5254gat = ~new_G5127gat & ~new_G5188gat;
  assign new_G5255gat = ~new_G5188gat & ~new_G723gat;
  assign new_G5256gat = ~new_G5017gat & ~new_G5188gat;
  assign new_G5259gat = ~new_G5192gat & ~new_G5193gat;
  assign new_G5262gat = ~new_G5197gat & ~new_G5194gat;
  assign new_G5266gat = ~new_G5139gat & ~new_G5200gat;
  assign new_G5267gat = ~new_G5200gat & ~new_G5136gat;
  assign new_G5268gat = ~new_G5204gat & ~new_G5205gat;
  assign new_G5271gat = ~new_G5206gat & ~new_G918gat;
  assign new_G5275gat = ~new_G5148gat & ~new_G5209gat;
  assign new_G5276gat = ~new_G5209gat & ~new_G966gat;
  assign new_G5277gat = ~new_G5038gat & ~new_G5209gat;
  assign new_G5280gat = ~new_G5213gat & ~new_G5214gat;
  assign new_G5283gat = ~new_G5218gat & ~new_G5215gat;
  assign new_G5287gat = ~new_G5160gat & ~new_G5221gat;
  assign new_G5288gat = ~new_G5221gat & ~new_G5157gat;
  assign new_G5289gat = ~new_G5225gat & ~new_G5226gat;
  assign new_G5292gat = ~new_G5227gat & ~new_G1161gat;
  assign new_G5296gat = ~new_G5169gat & ~new_G5230gat;
  assign new_G5297gat = ~new_G5230gat & ~new_G1209gat;
  assign new_G5298gat = ~new_G5059gat & ~new_G5230gat;
  assign new_G5301gat = ~new_G5234gat & ~new_G5235gat;
  assign new_G5304gat = ~new_G1305gat & ~new_G5236gat;
  assign G5308gat = ~new_G5239gat & ~new_G5240gat;
  assign new_G5309gat = ~new_G5244gat & ~new_G5245gat;
  assign new_G5312gat = ~new_G5249gat & ~new_G5250gat;
  assign new_G5315gat = ~new_G5254gat & ~new_G5255gat;
  assign new_G5318gat = ~new_G5259gat & ~new_G5256gat;
  assign new_G5322gat = ~new_G5197gat & ~new_G5262gat;
  assign new_G5323gat = ~new_G5262gat & ~new_G5194gat;
  assign new_G5324gat = ~new_G5266gat & ~new_G5267gat;
  assign new_G5327gat = ~new_G5268gat & ~new_G870gat;
  assign new_G5331gat = ~new_G5206gat & ~new_G5271gat;
  assign new_G5332gat = ~new_G5271gat & ~new_G918gat;
  assign new_G5333gat = ~new_G5088gat & ~new_G5271gat;
  assign new_G5336gat = ~new_G5275gat & ~new_G5276gat;
  assign new_G5339gat = ~new_G5280gat & ~new_G5277gat;
  assign new_G5343gat = ~new_G5218gat & ~new_G5283gat;
  assign new_G5344gat = ~new_G5283gat & ~new_G5215gat;
  assign new_G5345gat = ~new_G5287gat & ~new_G5288gat;
  assign new_G5348gat = ~new_G5289gat & ~new_G1113gat;
  assign new_G5352gat = ~new_G5227gat & ~new_G5292gat;
  assign new_G5353gat = ~new_G5292gat & ~new_G1161gat;
  assign new_G5354gat = ~new_G5109gat & ~new_G5292gat;
  assign new_G5357gat = ~new_G5296gat & ~new_G5297gat;
  assign new_G5360gat = ~new_G5301gat & ~new_G5298gat;
  assign new_G5364gat = ~new_G1305gat & ~new_G5304gat;
  assign new_G5365gat = ~new_G5304gat & ~new_G5236gat;
  assign new_G5366gat = ~new_G5309gat & ~new_G5241gat;
  assign new_G5370gat = ~new_G5312gat & ~new_G5246gat;
  assign new_G5374gat = ~new_G5315gat & ~new_G5251gat;
  assign new_G5378gat = ~new_G5259gat & ~new_G5318gat;
  assign new_G5379gat = ~new_G5318gat & ~new_G5256gat;
  assign new_G5380gat = ~new_G5322gat & ~new_G5323gat;
  assign new_G5383gat = ~new_G5324gat & ~new_G822gat;
  assign new_G5387gat = ~new_G5268gat & ~new_G5327gat;
  assign new_G5388gat = ~new_G5327gat & ~new_G870gat;
  assign new_G5389gat = ~new_G5142gat & ~new_G5327gat;
  assign new_G5392gat = ~new_G5331gat & ~new_G5332gat;
  assign new_G5395gat = ~new_G5336gat & ~new_G5333gat;
  assign new_G5399gat = ~new_G5280gat & ~new_G5339gat;
  assign new_G5400gat = ~new_G5339gat & ~new_G5277gat;
  assign new_G5401gat = ~new_G5343gat & ~new_G5344gat;
  assign new_G5404gat = ~new_G5345gat & ~new_G1065gat;
  assign new_G5408gat = ~new_G5289gat & ~new_G5348gat;
  assign new_G5409gat = ~new_G5348gat & ~new_G1113gat;
  assign new_G5410gat = ~new_G5163gat & ~new_G5348gat;
  assign new_G5413gat = ~new_G5352gat & ~new_G5353gat;
  assign new_G5416gat = ~new_G5357gat & ~new_G5354gat;
  assign new_G5420gat = ~new_G5301gat & ~new_G5360gat;
  assign new_G5421gat = ~new_G5360gat & ~new_G5298gat;
  assign new_G5422gat = ~new_G5364gat & ~new_G5365gat;
  assign new_G5425gat = ~new_G5309gat & ~new_G5366gat;
  assign new_G5426gat = ~new_G5366gat & ~new_G5241gat;
  assign new_G5427gat = ~new_G5312gat & ~new_G5370gat;
  assign new_G5428gat = ~new_G5370gat & ~new_G5246gat;
  assign new_G5429gat = ~new_G5315gat & ~new_G5374gat;
  assign new_G5430gat = ~new_G5374gat & ~new_G5251gat;
  assign new_G5431gat = ~new_G5378gat & ~new_G5379gat;
  assign new_G5434gat = ~new_G5380gat & ~new_G774gat;
  assign new_G5438gat = ~new_G5324gat & ~new_G5383gat;
  assign new_G5439gat = ~new_G5383gat & ~new_G822gat;
  assign new_G5440gat = ~new_G5200gat & ~new_G5383gat;
  assign new_G5443gat = ~new_G5387gat & ~new_G5388gat;
  assign new_G5446gat = ~new_G5392gat & ~new_G5389gat;
  assign new_G5450gat = ~new_G5336gat & ~new_G5395gat;
  assign new_G5451gat = ~new_G5395gat & ~new_G5333gat;
  assign new_G5452gat = ~new_G5399gat & ~new_G5400gat;
  assign new_G5455gat = ~new_G5401gat & ~new_G1017gat;
  assign new_G5459gat = ~new_G5345gat & ~new_G5404gat;
  assign new_G5460gat = ~new_G5404gat & ~new_G1065gat;
  assign new_G5461gat = ~new_G5221gat & ~new_G5404gat;
  assign new_G5464gat = ~new_G5408gat & ~new_G5409gat;
  assign new_G5467gat = ~new_G5413gat & ~new_G5410gat;
  assign new_G5471gat = ~new_G5357gat & ~new_G5416gat;
  assign new_G5472gat = ~new_G5416gat & ~new_G5354gat;
  assign new_G5473gat = ~new_G5420gat & ~new_G5421gat;
  assign new_G5476gat = ~new_G5422gat & ~new_G1260gat;
  assign new_G5480gat = ~new_G5425gat & ~new_G5426gat;
  assign new_G5483gat = ~new_G5427gat & ~new_G5428gat;
  assign new_G5486gat = ~new_G5429gat & ~new_G5430gat;
  assign new_G5489gat = ~new_G5431gat & ~new_G726gat;
  assign new_G5493gat = ~new_G5380gat & ~new_G5434gat;
  assign new_G5494gat = ~new_G5434gat & ~new_G774gat;
  assign new_G5495gat = ~new_G5262gat & ~new_G5434gat;
  assign new_G5498gat = ~new_G5438gat & ~new_G5439gat;
  assign new_G5501gat = ~new_G5443gat & ~new_G5440gat;
  assign new_G5505gat = ~new_G5392gat & ~new_G5446gat;
  assign new_G5506gat = ~new_G5446gat & ~new_G5389gat;
  assign new_G5507gat = ~new_G5450gat & ~new_G5451gat;
  assign new_G5510gat = ~new_G5452gat & ~new_G969gat;
  assign new_G5514gat = ~new_G5401gat & ~new_G5455gat;
  assign new_G5515gat = ~new_G5455gat & ~new_G1017gat;
  assign new_G5516gat = ~new_G5283gat & ~new_G5455gat;
  assign new_G5519gat = ~new_G5459gat & ~new_G5460gat;
  assign new_G5522gat = ~new_G5464gat & ~new_G5461gat;
  assign new_G5526gat = ~new_G5413gat & ~new_G5467gat;
  assign new_G5527gat = ~new_G5467gat & ~new_G5410gat;
  assign new_G5528gat = ~new_G5471gat & ~new_G5472gat;
  assign new_G5531gat = ~new_G5473gat & ~new_G1212gat;
  assign new_G5535gat = ~new_G5422gat & ~new_G5476gat;
  assign new_G5536gat = ~new_G5476gat & ~new_G1260gat;
  assign new_G5537gat = ~new_G5304gat & ~new_G5476gat;
  assign new_G5540gat = ~new_G5480gat & ~new_G582gat;
  assign new_G5544gat = ~new_G5483gat & ~new_G630gat;
  assign new_G5548gat = ~new_G5486gat & ~new_G678gat;
  assign new_G5552gat = ~new_G5431gat & ~new_G5489gat;
  assign new_G5553gat = ~new_G5489gat & ~new_G726gat;
  assign new_G5554gat = ~new_G5318gat & ~new_G5489gat;
  assign new_G5557gat = ~new_G5493gat & ~new_G5494gat;
  assign new_G5560gat = ~new_G5498gat & ~new_G5495gat;
  assign new_G5564gat = ~new_G5443gat & ~new_G5501gat;
  assign new_G5565gat = ~new_G5501gat & ~new_G5440gat;
  assign new_G5566gat = ~new_G5505gat & ~new_G5506gat;
  assign new_G5569gat = ~new_G5507gat & ~new_G921gat;
  assign new_G5573gat = ~new_G5452gat & ~new_G5510gat;
  assign new_G5574gat = ~new_G5510gat & ~new_G969gat;
  assign new_G5575gat = ~new_G5339gat & ~new_G5510gat;
  assign new_G5578gat = ~new_G5514gat & ~new_G5515gat;
  assign new_G5581gat = ~new_G5519gat & ~new_G5516gat;
  assign new_G5585gat = ~new_G5464gat & ~new_G5522gat;
  assign new_G5586gat = ~new_G5522gat & ~new_G5461gat;
  assign new_G5587gat = ~new_G5526gat & ~new_G5527gat;
  assign new_G5590gat = ~new_G5528gat & ~new_G1164gat;
  assign new_G5594gat = ~new_G5473gat & ~new_G5531gat;
  assign new_G5595gat = ~new_G5531gat & ~new_G1212gat;
  assign new_G5596gat = ~new_G5360gat & ~new_G5531gat;
  assign new_G5599gat = ~new_G5535gat & ~new_G5536gat;
  assign new_G5602gat = ~new_G1308gat & ~new_G5537gat;
  assign new_G5606gat = ~new_G5480gat & ~new_G5540gat;
  assign new_G5607gat = ~new_G5540gat & ~new_G582gat;
  assign new_G5608gat = ~new_G5366gat & ~new_G5540gat;
  assign new_G5611gat = ~new_G5483gat & ~new_G5544gat;
  assign new_G5612gat = ~new_G5544gat & ~new_G630gat;
  assign new_G5613gat = ~new_G5370gat & ~new_G5544gat;
  assign new_G5616gat = ~new_G5486gat & ~new_G5548gat;
  assign new_G5617gat = ~new_G5548gat & ~new_G678gat;
  assign new_G5618gat = ~new_G5374gat & ~new_G5548gat;
  assign new_G5621gat = ~new_G5552gat & ~new_G5553gat;
  assign new_G5624gat = ~new_G5557gat & ~new_G5554gat;
  assign new_G5628gat = ~new_G5498gat & ~new_G5560gat;
  assign new_G5629gat = ~new_G5560gat & ~new_G5495gat;
  assign new_G5630gat = ~new_G5564gat & ~new_G5565gat;
  assign new_G5633gat = ~new_G5566gat & ~new_G873gat;
  assign new_G5637gat = ~new_G5507gat & ~new_G5569gat;
  assign new_G5638gat = ~new_G5569gat & ~new_G921gat;
  assign new_G5639gat = ~new_G5395gat & ~new_G5569gat;
  assign new_G5642gat = ~new_G5573gat & ~new_G5574gat;
  assign new_G5645gat = ~new_G5578gat & ~new_G5575gat;
  assign new_G5649gat = ~new_G5519gat & ~new_G5581gat;
  assign new_G5650gat = ~new_G5581gat & ~new_G5516gat;
  assign new_G5651gat = ~new_G5585gat & ~new_G5586gat;
  assign new_G5654gat = ~new_G5587gat & ~new_G1116gat;
  assign new_G5658gat = ~new_G5528gat & ~new_G5590gat;
  assign new_G5659gat = ~new_G5590gat & ~new_G1164gat;
  assign new_G5660gat = ~new_G5416gat & ~new_G5590gat;
  assign new_G5663gat = ~new_G5594gat & ~new_G5595gat;
  assign new_G5666gat = ~new_G5599gat & ~new_G5596gat;
  assign new_G5670gat = ~new_G1308gat & ~new_G5602gat;
  assign new_G5671gat = ~new_G5602gat & ~new_G5537gat;
  assign G5672gat = ~new_G5606gat & ~new_G5607gat;
  assign new_G5673gat = ~new_G5611gat & ~new_G5612gat;
  assign new_G5676gat = ~new_G5616gat & ~new_G5617gat;
  assign new_G5679gat = ~new_G5621gat & ~new_G5618gat;
  assign new_G5683gat = ~new_G5557gat & ~new_G5624gat;
  assign new_G5684gat = ~new_G5624gat & ~new_G5554gat;
  assign new_G5685gat = ~new_G5628gat & ~new_G5629gat;
  assign new_G5688gat = ~new_G5630gat & ~new_G825gat;
  assign new_G5692gat = ~new_G5566gat & ~new_G5633gat;
  assign new_G5693gat = ~new_G5633gat & ~new_G873gat;
  assign new_G5694gat = ~new_G5446gat & ~new_G5633gat;
  assign new_G5697gat = ~new_G5637gat & ~new_G5638gat;
  assign new_G5700gat = ~new_G5642gat & ~new_G5639gat;
  assign new_G5704gat = ~new_G5578gat & ~new_G5645gat;
  assign new_G5705gat = ~new_G5645gat & ~new_G5575gat;
  assign new_G5706gat = ~new_G5649gat & ~new_G5650gat;
  assign new_G5709gat = ~new_G5651gat & ~new_G1068gat;
  assign new_G5713gat = ~new_G5587gat & ~new_G5654gat;
  assign new_G5714gat = ~new_G5654gat & ~new_G1116gat;
  assign new_G5715gat = ~new_G5467gat & ~new_G5654gat;
  assign new_G5718gat = ~new_G5658gat & ~new_G5659gat;
  assign new_G5721gat = ~new_G5663gat & ~new_G5660gat;
  assign new_G5725gat = ~new_G5599gat & ~new_G5666gat;
  assign new_G5726gat = ~new_G5666gat & ~new_G5596gat;
  assign new_G5727gat = ~new_G5670gat & ~new_G5671gat;
  assign new_G5730gat = ~new_G5673gat & ~new_G5608gat;
  assign new_G5734gat = ~new_G5676gat & ~new_G5613gat;
  assign new_G5738gat = ~new_G5621gat & ~new_G5679gat;
  assign new_G5739gat = ~new_G5679gat & ~new_G5618gat;
  assign new_G5740gat = ~new_G5683gat & ~new_G5684gat;
  assign new_G5743gat = ~new_G5685gat & ~new_G777gat;
  assign new_G5747gat = ~new_G5630gat & ~new_G5688gat;
  assign new_G5748gat = ~new_G5688gat & ~new_G825gat;
  assign new_G5749gat = ~new_G5501gat & ~new_G5688gat;
  assign new_G5752gat = ~new_G5692gat & ~new_G5693gat;
  assign new_G5755gat = ~new_G5697gat & ~new_G5694gat;
  assign new_G5759gat = ~new_G5642gat & ~new_G5700gat;
  assign new_G5760gat = ~new_G5700gat & ~new_G5639gat;
  assign new_G5761gat = ~new_G5704gat & ~new_G5705gat;
  assign new_G5764gat = ~new_G5706gat & ~new_G1020gat;
  assign new_G5768gat = ~new_G5651gat & ~new_G5709gat;
  assign new_G5769gat = ~new_G5709gat & ~new_G1068gat;
  assign new_G5770gat = ~new_G5522gat & ~new_G5709gat;
  assign new_G5773gat = ~new_G5713gat & ~new_G5714gat;
  assign new_G5776gat = ~new_G5718gat & ~new_G5715gat;
  assign new_G5780gat = ~new_G5663gat & ~new_G5721gat;
  assign new_G5781gat = ~new_G5721gat & ~new_G5660gat;
  assign new_G5782gat = ~new_G5725gat & ~new_G5726gat;
  assign new_G5785gat = ~new_G5673gat & ~new_G5730gat;
  assign new_G5786gat = ~new_G5730gat & ~new_G5608gat;
  assign new_G5787gat = ~new_G5676gat & ~new_G5734gat;
  assign new_G5788gat = ~new_G5734gat & ~new_G5613gat;
  assign new_G5789gat = ~new_G5738gat & ~new_G5739gat;
  assign new_G5792gat = ~new_G5740gat & ~new_G729gat;
  assign new_G5796gat = ~new_G5685gat & ~new_G5743gat;
  assign new_G5797gat = ~new_G5743gat & ~new_G777gat;
  assign new_G5798gat = ~new_G5560gat & ~new_G5743gat;
  assign new_G5801gat = ~new_G5747gat & ~new_G5748gat;
  assign new_G5804gat = ~new_G5752gat & ~new_G5749gat;
  assign new_G5808gat = ~new_G5697gat & ~new_G5755gat;
  assign new_G5809gat = ~new_G5755gat & ~new_G5694gat;
  assign new_G5810gat = ~new_G5759gat & ~new_G5760gat;
  assign new_G5813gat = ~new_G5761gat & ~new_G972gat;
  assign new_G5817gat = ~new_G5706gat & ~new_G5764gat;
  assign new_G5818gat = ~new_G5764gat & ~new_G1020gat;
  assign new_G5819gat = ~new_G5581gat & ~new_G5764gat;
  assign new_G5822gat = ~new_G5768gat & ~new_G5769gat;
  assign new_G5825gat = ~new_G5773gat & ~new_G5770gat;
  assign new_G5829gat = ~new_G5718gat & ~new_G5776gat;
  assign new_G5830gat = ~new_G5776gat & ~new_G5715gat;
  assign new_G5831gat = ~new_G5780gat & ~new_G5781gat;
  assign new_G5834gat = ~new_G5785gat & ~new_G5786gat;
  assign new_G5837gat = ~new_G5787gat & ~new_G5788gat;
  assign new_G5840gat = ~new_G5789gat & ~new_G681gat;
  assign new_G5844gat = ~new_G5740gat & ~new_G5792gat;
  assign new_G5845gat = ~new_G5792gat & ~new_G729gat;
  assign new_G5846gat = ~new_G5624gat & ~new_G5792gat;
  assign new_G5849gat = ~new_G5796gat & ~new_G5797gat;
  assign new_G5852gat = ~new_G5801gat & ~new_G5798gat;
  assign new_G5856gat = ~new_G5752gat & ~new_G5804gat;
  assign new_G5857gat = ~new_G5804gat & ~new_G5749gat;
  assign new_G5858gat = ~new_G5808gat & ~new_G5809gat;
  assign new_G5861gat = ~new_G5810gat & ~new_G924gat;
  assign new_G5865gat = ~new_G5761gat & ~new_G5813gat;
  assign new_G5866gat = ~new_G5813gat & ~new_G972gat;
  assign new_G5867gat = ~new_G5645gat & ~new_G5813gat;
  assign new_G5870gat = ~new_G5817gat & ~new_G5818gat;
  assign new_G5873gat = ~new_G5822gat & ~new_G5819gat;
  assign new_G5877gat = ~new_G5773gat & ~new_G5825gat;
  assign new_G5878gat = ~new_G5825gat & ~new_G5770gat;
  assign new_G5879gat = ~new_G5829gat & ~new_G5830gat;
  assign new_G5882gat = ~new_G5834gat & ~new_G585gat;
  assign new_G5886gat = ~new_G5837gat & ~new_G633gat;
  assign new_G5890gat = ~new_G5789gat & ~new_G5840gat;
  assign new_G5891gat = ~new_G5840gat & ~new_G681gat;
  assign new_G5892gat = ~new_G5679gat & ~new_G5840gat;
  assign new_G5895gat = ~new_G5844gat & ~new_G5845gat;
  assign new_G5898gat = ~new_G5849gat & ~new_G5846gat;
  assign new_G5902gat = ~new_G5801gat & ~new_G5852gat;
  assign new_G5903gat = ~new_G5852gat & ~new_G5798gat;
  assign new_G5904gat = ~new_G5856gat & ~new_G5857gat;
  assign new_G5907gat = ~new_G5858gat & ~new_G876gat;
  assign new_G5911gat = ~new_G5810gat & ~new_G5861gat;
  assign new_G5912gat = ~new_G5861gat & ~new_G924gat;
  assign new_G5913gat = ~new_G5700gat & ~new_G5861gat;
  assign new_G5916gat = ~new_G5865gat & ~new_G5866gat;
  assign new_G5919gat = ~new_G5870gat & ~new_G5867gat;
  assign new_G5923gat = ~new_G5822gat & ~new_G5873gat;
  assign new_G5924gat = ~new_G5873gat & ~new_G5819gat;
  assign new_G5925gat = ~new_G5877gat & ~new_G5878gat;
  assign new_G5928gat = ~new_G5834gat & ~new_G5882gat;
  assign new_G5929gat = ~new_G5882gat & ~new_G585gat;
  assign new_G5930gat = ~new_G5730gat & ~new_G5882gat;
  assign new_G5933gat = ~new_G5837gat & ~new_G5886gat;
  assign new_G5934gat = ~new_G5886gat & ~new_G633gat;
  assign new_G5935gat = ~new_G5734gat & ~new_G5886gat;
  assign new_G5938gat = ~new_G5890gat & ~new_G5891gat;
  assign new_G5941gat = ~new_G5895gat & ~new_G5892gat;
  assign new_G5945gat = ~new_G5849gat & ~new_G5898gat;
  assign new_G5946gat = ~new_G5898gat & ~new_G5846gat;
  assign new_G5947gat = ~new_G5902gat & ~new_G5903gat;
  assign new_G5950gat = ~new_G5904gat & ~new_G828gat;
  assign new_G5954gat = ~new_G5858gat & ~new_G5907gat;
  assign new_G5955gat = ~new_G5907gat & ~new_G876gat;
  assign new_G5956gat = ~new_G5755gat & ~new_G5907gat;
  assign new_G5959gat = ~new_G5911gat & ~new_G5912gat;
  assign new_G5962gat = ~new_G5916gat & ~new_G5913gat;
  assign new_G5966gat = ~new_G5870gat & ~new_G5919gat;
  assign new_G5967gat = ~new_G5919gat & ~new_G5867gat;
  assign new_G5968gat = ~new_G5923gat & ~new_G5924gat;
  assign G5971gat = ~new_G5928gat & ~new_G5929gat;
  assign new_G5972gat = ~new_G5933gat & ~new_G5934gat;
  assign new_G5975gat = ~new_G5938gat & ~new_G5935gat;
  assign new_G5979gat = ~new_G5895gat & ~new_G5941gat;
  assign new_G5980gat = ~new_G5941gat & ~new_G5892gat;
  assign new_G5981gat = ~new_G5945gat & ~new_G5946gat;
  assign new_G5984gat = ~new_G5947gat & ~new_G780gat;
  assign new_G5988gat = ~new_G5904gat & ~new_G5950gat;
  assign new_G5989gat = ~new_G5950gat & ~new_G828gat;
  assign new_G5990gat = ~new_G5804gat & ~new_G5950gat;
  assign new_G5993gat = ~new_G5954gat & ~new_G5955gat;
  assign new_G5996gat = ~new_G5959gat & ~new_G5956gat;
  assign new_G6000gat = ~new_G5916gat & ~new_G5962gat;
  assign new_G6001gat = ~new_G5962gat & ~new_G5913gat;
  assign new_G6002gat = ~new_G5966gat & ~new_G5967gat;
  assign new_G6005gat = ~new_G5972gat & ~new_G5930gat;
  assign new_G6009gat = ~new_G5938gat & ~new_G5975gat;
  assign new_G6010gat = ~new_G5975gat & ~new_G5935gat;
  assign new_G6011gat = ~new_G5979gat & ~new_G5980gat;
  assign new_G6014gat = ~new_G5981gat & ~new_G732gat;
  assign new_G6018gat = ~new_G5947gat & ~new_G5984gat;
  assign new_G6019gat = ~new_G5984gat & ~new_G780gat;
  assign new_G6020gat = ~new_G5852gat & ~new_G5984gat;
  assign new_G6023gat = ~new_G5988gat & ~new_G5989gat;
  assign new_G6026gat = ~new_G5993gat & ~new_G5990gat;
  assign new_G6030gat = ~new_G5959gat & ~new_G5996gat;
  assign new_G6031gat = ~new_G5996gat & ~new_G5956gat;
  assign new_G6032gat = ~new_G6000gat & ~new_G6001gat;
  assign new_G6035gat = ~new_G5972gat & ~new_G6005gat;
  assign new_G6036gat = ~new_G6005gat & ~new_G5930gat;
  assign new_G6037gat = ~new_G6009gat & ~new_G6010gat;
  assign new_G6040gat = ~new_G6011gat & ~new_G684gat;
  assign new_G6044gat = ~new_G5981gat & ~new_G6014gat;
  assign new_G6045gat = ~new_G6014gat & ~new_G732gat;
  assign new_G6046gat = ~new_G5898gat & ~new_G6014gat;
  assign new_G6049gat = ~new_G6018gat & ~new_G6019gat;
  assign new_G6052gat = ~new_G6023gat & ~new_G6020gat;
  assign new_G6056gat = ~new_G5993gat & ~new_G6026gat;
  assign new_G6057gat = ~new_G6026gat & ~new_G5990gat;
  assign new_G6058gat = ~new_G6030gat & ~new_G6031gat;
  assign new_G6061gat = ~new_G6035gat & ~new_G6036gat;
  assign new_G6064gat = ~new_G6037gat & ~new_G636gat;
  assign new_G6068gat = ~new_G6011gat & ~new_G6040gat;
  assign new_G6069gat = ~new_G6040gat & ~new_G684gat;
  assign new_G6070gat = ~new_G5941gat & ~new_G6040gat;
  assign new_G6073gat = ~new_G6044gat & ~new_G6045gat;
  assign new_G6076gat = ~new_G6049gat & ~new_G6046gat;
  assign new_G6080gat = ~new_G6023gat & ~new_G6052gat;
  assign new_G6081gat = ~new_G6052gat & ~new_G6020gat;
  assign new_G6082gat = ~new_G6056gat & ~new_G6057gat;
  assign new_G6085gat = ~new_G6061gat & ~new_G588gat;
  assign new_G6089gat = ~new_G6037gat & ~new_G6064gat;
  assign new_G6090gat = ~new_G6064gat & ~new_G636gat;
  assign new_G6091gat = ~new_G5975gat & ~new_G6064gat;
  assign new_G6094gat = ~new_G6068gat & ~new_G6069gat;
  assign new_G6097gat = ~new_G6073gat & ~new_G6070gat;
  assign new_G6101gat = ~new_G6049gat & ~new_G6076gat;
  assign new_G6102gat = ~new_G6076gat & ~new_G6046gat;
  assign new_G6103gat = ~new_G6080gat & ~new_G6081gat;
  assign new_G6106gat = ~new_G6061gat & ~new_G6085gat;
  assign new_G6107gat = ~new_G6085gat & ~new_G588gat;
  assign new_G6108gat = ~new_G6005gat & ~new_G6085gat;
  assign new_G6111gat = ~new_G6089gat & ~new_G6090gat;
  assign new_G6114gat = ~new_G6094gat & ~new_G6091gat;
  assign new_G6118gat = ~new_G6073gat & ~new_G6097gat;
  assign new_G6119gat = ~new_G6097gat & ~new_G6070gat;
  assign new_G6120gat = ~new_G6101gat & ~new_G6102gat;
  assign G6123gat = ~new_G6106gat & ~new_G6107gat;
  assign new_G6124gat = ~new_G6111gat & ~new_G6108gat;
  assign new_G6128gat = ~new_G6094gat & ~new_G6114gat;
  assign new_G6129gat = ~new_G6114gat & ~new_G6091gat;
  assign new_G6130gat = ~new_G6118gat & ~new_G6119gat;
  assign new_G6133gat = ~new_G6111gat & ~new_G6124gat;
  assign new_G6134gat = ~new_G6124gat & ~new_G6108gat;
  assign new_G6135gat = ~new_G6128gat & ~new_G6129gat;
  assign new_G6138gat = ~new_G6133gat & ~new_G6134gat;
  assign new_G6141gat = ~new_G6138gat;
  assign new_G6145gat = ~new_G6138gat & ~new_G6141gat;
  assign new_G6146gat = ~new_G6141gat;
  assign new_G6147gat = ~new_G6124gat & ~new_G6141gat;
  assign G6150gat = ~new_G6145gat & ~new_G6146gat;
  assign new_G6151gat = ~new_G6135gat & ~new_G6147gat;
  assign new_G6155gat = ~new_G6135gat & ~new_G6151gat;
  assign new_G6156gat = ~new_G6151gat & ~new_G6147gat;
  assign new_G6157gat = ~new_G6114gat & ~new_G6151gat;
  assign G6160gat = ~new_G6155gat & ~new_G6156gat;
  assign new_G6161gat = ~new_G6130gat & ~new_G6157gat;
  assign new_G6165gat = ~new_G6130gat & ~new_G6161gat;
  assign new_G6166gat = ~new_G6161gat & ~new_G6157gat;
  assign new_G6167gat = ~new_G6097gat & ~new_G6161gat;
  assign G6170gat = ~new_G6165gat & ~new_G6166gat;
  assign new_G6171gat = ~new_G6120gat & ~new_G6167gat;
  assign new_G6175gat = ~new_G6120gat & ~new_G6171gat;
  assign new_G6176gat = ~new_G6171gat & ~new_G6167gat;
  assign new_G6177gat = ~new_G6076gat & ~new_G6171gat;
  assign G6180gat = ~new_G6175gat & ~new_G6176gat;
  assign new_G6181gat = ~new_G6103gat & ~new_G6177gat;
  assign new_G6185gat = ~new_G6103gat & ~new_G6181gat;
  assign new_G6186gat = ~new_G6181gat & ~new_G6177gat;
  assign new_G6187gat = ~new_G6052gat & ~new_G6181gat;
  assign G6190gat = ~new_G6185gat & ~new_G6186gat;
  assign new_G6191gat = ~new_G6082gat & ~new_G6187gat;
  assign new_G6195gat = ~new_G6082gat & ~new_G6191gat;
  assign new_G6196gat = ~new_G6191gat & ~new_G6187gat;
  assign new_G6197gat = ~new_G6026gat & ~new_G6191gat;
  assign G6200gat = ~new_G6195gat & ~new_G6196gat;
  assign new_G6201gat = ~new_G6058gat & ~new_G6197gat;
  assign new_G6205gat = ~new_G6058gat & ~new_G6201gat;
  assign new_G6206gat = ~new_G6201gat & ~new_G6197gat;
  assign new_G6207gat = ~new_G5996gat & ~new_G6201gat;
  assign G6210gat = ~new_G6205gat & ~new_G6206gat;
  assign new_G6211gat = ~new_G6032gat & ~new_G6207gat;
  assign new_G6215gat = ~new_G6032gat & ~new_G6211gat;
  assign new_G6216gat = ~new_G6211gat & ~new_G6207gat;
  assign new_G6217gat = ~new_G5962gat & ~new_G6211gat;
  assign G6220gat = ~new_G6215gat & ~new_G6216gat;
  assign new_G6221gat = ~new_G6002gat & ~new_G6217gat;
  assign new_G6225gat = ~new_G6002gat & ~new_G6221gat;
  assign new_G6226gat = ~new_G6221gat & ~new_G6217gat;
  assign new_G6227gat = ~new_G5919gat & ~new_G6221gat;
  assign G6230gat = ~new_G6225gat & ~new_G6226gat;
  assign new_G6231gat = ~new_G5968gat & ~new_G6227gat;
  assign new_G6235gat = ~new_G5968gat & ~new_G6231gat;
  assign new_G6236gat = ~new_G6231gat & ~new_G6227gat;
  assign new_G6237gat = ~new_G5873gat & ~new_G6231gat;
  assign G6240gat = ~new_G6235gat & ~new_G6236gat;
  assign new_G6241gat = ~new_G5925gat & ~new_G6237gat;
  assign new_G6245gat = ~new_G5925gat & ~new_G6241gat;
  assign new_G6246gat = ~new_G6241gat & ~new_G6237gat;
  assign new_G6247gat = ~new_G5825gat & ~new_G6241gat;
  assign G6250gat = ~new_G6245gat & ~new_G6246gat;
  assign new_G6251gat = ~new_G5879gat & ~new_G6247gat;
  assign new_G6255gat = ~new_G5879gat & ~new_G6251gat;
  assign new_G6256gat = ~new_G6251gat & ~new_G6247gat;
  assign new_G6257gat = ~new_G5776gat & ~new_G6251gat;
  assign G6260gat = ~new_G6255gat & ~new_G6256gat;
  assign new_G6261gat = ~new_G5831gat & ~new_G6257gat;
  assign new_G6265gat = ~new_G5831gat & ~new_G6261gat;
  assign new_G6266gat = ~new_G6261gat & ~new_G6257gat;
  assign new_G6267gat = ~new_G5721gat & ~new_G6261gat;
  assign G6270gat = ~new_G6265gat & ~new_G6266gat;
  assign new_G6271gat = ~new_G5782gat & ~new_G6267gat;
  assign new_G6275gat = ~new_G5782gat & ~new_G6271gat;
  assign new_G6276gat = ~new_G6271gat & ~new_G6267gat;
  assign new_G6277gat = ~new_G5666gat & ~new_G6271gat;
  assign G6280gat = ~new_G6275gat & ~new_G6276gat;
  assign new_G6281gat = ~new_G5727gat & ~new_G6277gat;
  assign new_G6285gat = ~new_G5727gat & ~new_G6281gat;
  assign new_G6286gat = ~new_G6281gat & ~new_G6277gat;
  assign G6287gat = ~new_G5602gat & ~new_G6281gat;
  assign G6288gat = ~new_G6285gat & ~new_G6286gat;
endmodule
