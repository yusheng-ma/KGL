// Benchmark "./benchmarks/iscas85/c1355" written by ABC on Sun Apr 28 12:32:37 2024

module c1355  ( 
    G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
    G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
    G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat,
    G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat,
    G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat,
    G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat,
    G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
    G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat,
    G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat,
    G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_G242gat, new_G245gat, new_G248gat, new_G251gat, new_G254gat,
    new_G257gat, new_G260gat, new_G263gat, new_G266gat, new_G269gat,
    new_G272gat, new_G275gat, new_G278gat, new_G281gat, new_G284gat,
    new_G287gat, new_G290gat, new_G293gat, new_G296gat, new_G299gat,
    new_G302gat, new_G305gat, new_G308gat, new_G311gat, new_G314gat,
    new_G317gat, new_G320gat, new_G323gat, new_G326gat, new_G329gat,
    new_G332gat, new_G335gat, new_G338gat, new_G341gat, new_G344gat,
    new_G347gat, new_G350gat, new_G353gat, new_G356gat, new_G359gat,
    new_G362gat, new_G363gat, new_G364gat, new_G365gat, new_G366gat,
    new_G367gat, new_G368gat, new_G369gat, new_G370gat, new_G371gat,
    new_G372gat, new_G373gat, new_G374gat, new_G375gat, new_G376gat,
    new_G377gat, new_G378gat, new_G379gat, new_G380gat, new_G381gat,
    new_G382gat, new_G383gat, new_G384gat, new_G385gat, new_G386gat,
    new_G387gat, new_G388gat, new_G389gat, new_G390gat, new_G391gat,
    new_G392gat, new_G393gat, new_G394gat, new_G395gat, new_G396gat,
    new_G397gat, new_G398gat, new_G399gat, new_G400gat, new_G401gat,
    new_G402gat, new_G403gat, new_G404gat, new_G405gat, new_G406gat,
    new_G407gat, new_G408gat, new_G409gat, new_G410gat, new_G411gat,
    new_G412gat, new_G413gat, new_G414gat, new_G415gat, new_G416gat,
    new_G417gat, new_G418gat, new_G419gat, new_G420gat, new_G421gat,
    new_G422gat, new_G423gat, new_G424gat, new_G425gat, new_G426gat,
    new_G429gat, new_G432gat, new_G435gat, new_G438gat, new_G441gat,
    new_G444gat, new_G447gat, new_G450gat, new_G453gat, new_G456gat,
    new_G459gat, new_G462gat, new_G465gat, new_G468gat, new_G471gat,
    new_G474gat, new_G477gat, new_G480gat, new_G483gat, new_G486gat,
    new_G489gat, new_G492gat, new_G495gat, new_G498gat, new_G501gat,
    new_G504gat, new_G507gat, new_G510gat, new_G513gat, new_G516gat,
    new_G519gat, new_G522gat, new_G525gat, new_G528gat, new_G531gat,
    new_G534gat, new_G537gat, new_G540gat, new_G543gat, new_G546gat,
    new_G549gat, new_G552gat, new_G555gat, new_G558gat, new_G561gat,
    new_G564gat, new_G567gat, new_G570gat, new_G571gat, new_G572gat,
    new_G573gat, new_G574gat, new_G575gat, new_G576gat, new_G577gat,
    new_G578gat, new_G579gat, new_G580gat, new_G581gat, new_G582gat,
    new_G583gat, new_G584gat, new_G585gat, new_G586gat, new_G587gat,
    new_G588gat, new_G589gat, new_G590gat, new_G591gat, new_G592gat,
    new_G593gat, new_G594gat, new_G595gat, new_G596gat, new_G597gat,
    new_G598gat, new_G599gat, new_G600gat, new_G601gat, new_G602gat,
    new_G607gat, new_G612gat, new_G617gat, new_G622gat, new_G627gat,
    new_G632gat, new_G637gat, new_G642gat, new_G645gat, new_G648gat,
    new_G651gat, new_G654gat, new_G657gat, new_G660gat, new_G663gat,
    new_G666gat, new_G669gat, new_G672gat, new_G675gat, new_G678gat,
    new_G681gat, new_G684gat, new_G687gat, new_G690gat, new_G691gat,
    new_G692gat, new_G693gat, new_G694gat, new_G695gat, new_G696gat,
    new_G697gat, new_G698gat, new_G699gat, new_G700gat, new_G701gat,
    new_G702gat, new_G703gat, new_G704gat, new_G705gat, new_G706gat,
    new_G709gat, new_G712gat, new_G715gat, new_G718gat, new_G721gat,
    new_G724gat, new_G727gat, new_G730gat, new_G733gat, new_G736gat,
    new_G739gat, new_G742gat, new_G745gat, new_G748gat, new_G751gat,
    new_G754gat, new_G755gat, new_G756gat, new_G757gat, new_G758gat,
    new_G759gat, new_G760gat, new_G761gat, new_G762gat, new_G763gat,
    new_G764gat, new_G765gat, new_G766gat, new_G767gat, new_G768gat,
    new_G769gat, new_G770gat, new_G773gat, new_G776gat, new_G779gat,
    new_G782gat, new_G785gat, new_G788gat, new_G791gat, new_G794gat,
    new_G797gat, new_G800gat, new_G803gat, new_G806gat, new_G809gat,
    new_G812gat, new_G815gat, new_G818gat, new_G819gat, new_G820gat,
    new_G821gat, new_G822gat, new_G823gat, new_G824gat, new_G825gat,
    new_G826gat, new_G827gat, new_G828gat, new_G829gat, new_G830gat,
    new_G831gat, new_G832gat, new_G833gat, new_G834gat, new_G847gat,
    new_G860gat, new_G873gat, new_G886gat, new_G899gat, new_G912gat,
    new_G925gat, new_G938gat, new_G939gat, new_G940gat, new_G941gat,
    new_G942gat, new_G943gat, new_G944gat, new_G945gat, new_G946gat,
    new_G947gat, new_G948gat, new_G949gat, new_G950gat, new_G951gat,
    new_G952gat, new_G953gat, new_G954gat, new_G955gat, new_G956gat,
    new_G957gat, new_G958gat, new_G959gat, new_G960gat, new_G961gat,
    new_G962gat, new_G963gat, new_G964gat, new_G965gat, new_G966gat,
    new_G967gat, new_G968gat, new_G969gat, new_G970gat, new_G971gat,
    new_G972gat, new_G973gat, new_G974gat, new_G975gat, new_G976gat,
    new_G977gat, new_G978gat, new_G979gat, new_G980gat, new_G981gat,
    new_G982gat, new_G983gat, new_G984gat, new_G985gat, new_G986gat,
    new_G991gat, new_G996gat, new_G1001gat, new_G1006gat, new_G1011gat,
    new_G1016gat, new_G1021gat, new_G1026gat, new_G1031gat, new_G1036gat,
    new_G1039gat, new_G1042gat, new_G1045gat, new_G1048gat, new_G1051gat,
    new_G1054gat, new_G1057gat, new_G1060gat, new_G1063gat, new_G1066gat,
    new_G1069gat, new_G1072gat, new_G1075gat, new_G1078gat, new_G1081gat,
    new_G1084gat, new_G1087gat, new_G1090gat, new_G1093gat, new_G1096gat,
    new_G1099gat, new_G1102gat, new_G1105gat, new_G1108gat, new_G1111gat,
    new_G1114gat, new_G1117gat, new_G1120gat, new_G1123gat, new_G1126gat,
    new_G1129gat, new_G1132gat, new_G1135gat, new_G1138gat, new_G1141gat,
    new_G1144gat, new_G1147gat, new_G1150gat, new_G1153gat, new_G1156gat,
    new_G1159gat, new_G1162gat, new_G1165gat, new_G1168gat, new_G1171gat,
    new_G1174gat, new_G1177gat, new_G1180gat, new_G1183gat, new_G1186gat,
    new_G1189gat, new_G1192gat, new_G1195gat, new_G1198gat, new_G1201gat,
    new_G1204gat, new_G1207gat, new_G1210gat, new_G1213gat, new_G1216gat,
    new_G1219gat, new_G1222gat, new_G1225gat, new_G1228gat, new_G1229gat,
    new_G1230gat, new_G1231gat, new_G1232gat, new_G1233gat, new_G1234gat,
    new_G1235gat, new_G1236gat, new_G1237gat, new_G1238gat, new_G1239gat,
    new_G1240gat, new_G1241gat, new_G1242gat, new_G1243gat, new_G1244gat,
    new_G1245gat, new_G1246gat, new_G1247gat, new_G1248gat, new_G1249gat,
    new_G1250gat, new_G1251gat, new_G1252gat, new_G1253gat, new_G1254gat,
    new_G1255gat, new_G1256gat, new_G1257gat, new_G1258gat, new_G1259gat,
    new_G1260gat, new_G1261gat, new_G1262gat, new_G1263gat, new_G1264gat,
    new_G1265gat, new_G1266gat, new_G1267gat, new_G1268gat, new_G1269gat,
    new_G1270gat, new_G1271gat, new_G1272gat, new_G1273gat, new_G1274gat,
    new_G1275gat, new_G1276gat, new_G1277gat, new_G1278gat, new_G1279gat,
    new_G1280gat, new_G1281gat, new_G1282gat, new_G1283gat, new_G1284gat,
    new_G1285gat, new_G1286gat, new_G1287gat, new_G1288gat, new_G1289gat,
    new_G1290gat, new_G1291gat, new_G1292gat, new_G1293gat, new_G1294gat,
    new_G1295gat, new_G1296gat, new_G1297gat, new_G1298gat, new_G1299gat,
    new_G1300gat, new_G1301gat, new_G1302gat, new_G1303gat, new_G1304gat,
    new_G1305gat, new_G1306gat, new_G1307gat, new_G1308gat, new_G1309gat,
    new_G1310gat, new_G1311gat, new_G1312gat, new_G1313gat, new_G1314gat,
    new_G1315gat, new_G1316gat, new_G1317gat, new_G1318gat, new_G1319gat,
    new_G1320gat, new_G1321gat, new_G1322gat, new_G1323gat;
  assign new_G242gat = G225gat & G233gat;
  assign new_G245gat = G226gat & G233gat;
  assign new_G248gat = G227gat & G233gat;
  assign new_G251gat = G228gat & G233gat;
  assign new_G254gat = G229gat & G233gat;
  assign new_G257gat = G230gat & G233gat;
  assign new_G260gat = G231gat & G233gat;
  assign new_G263gat = G232gat & G233gat;
  assign new_G266gat = ~G1gat | ~G8gat;
  assign new_G269gat = ~G15gat | ~G22gat;
  assign new_G272gat = ~G29gat | ~G36gat;
  assign new_G275gat = ~G43gat | ~G50gat;
  assign new_G278gat = ~G57gat | ~G64gat;
  assign new_G281gat = ~G71gat | ~G78gat;
  assign new_G284gat = ~G85gat | ~G92gat;
  assign new_G287gat = ~G99gat | ~G106gat;
  assign new_G290gat = ~G113gat | ~G120gat;
  assign new_G293gat = ~G127gat | ~G134gat;
  assign new_G296gat = ~G141gat | ~G148gat;
  assign new_G299gat = ~G155gat | ~G162gat;
  assign new_G302gat = ~G169gat | ~G176gat;
  assign new_G305gat = ~G183gat | ~G190gat;
  assign new_G308gat = ~G197gat | ~G204gat;
  assign new_G311gat = ~G211gat | ~G218gat;
  assign new_G314gat = ~G1gat | ~G29gat;
  assign new_G317gat = ~G57gat | ~G85gat;
  assign new_G320gat = ~G8gat | ~G36gat;
  assign new_G323gat = ~G64gat | ~G92gat;
  assign new_G326gat = ~G15gat | ~G43gat;
  assign new_G329gat = ~G71gat | ~G99gat;
  assign new_G332gat = ~G22gat | ~G50gat;
  assign new_G335gat = ~G78gat | ~G106gat;
  assign new_G338gat = ~G113gat | ~G141gat;
  assign new_G341gat = ~G169gat | ~G197gat;
  assign new_G344gat = ~G120gat | ~G148gat;
  assign new_G347gat = ~G176gat | ~G204gat;
  assign new_G350gat = ~G127gat | ~G155gat;
  assign new_G353gat = ~G183gat | ~G211gat;
  assign new_G356gat = ~G134gat | ~G162gat;
  assign new_G359gat = ~G190gat | ~G218gat;
  assign new_G362gat = ~G1gat | ~new_G266gat;
  assign new_G363gat = ~G8gat | ~new_G266gat;
  assign new_G364gat = ~G15gat | ~new_G269gat;
  assign new_G365gat = ~G22gat | ~new_G269gat;
  assign new_G366gat = ~G29gat | ~new_G272gat;
  assign new_G367gat = ~G36gat | ~new_G272gat;
  assign new_G368gat = ~G43gat | ~new_G275gat;
  assign new_G369gat = ~G50gat | ~new_G275gat;
  assign new_G370gat = ~G57gat | ~new_G278gat;
  assign new_G371gat = ~G64gat | ~new_G278gat;
  assign new_G372gat = ~G71gat | ~new_G281gat;
  assign new_G373gat = ~G78gat | ~new_G281gat;
  assign new_G374gat = ~G85gat | ~new_G284gat;
  assign new_G375gat = ~G92gat | ~new_G284gat;
  assign new_G376gat = ~G99gat | ~new_G287gat;
  assign new_G377gat = ~G106gat | ~new_G287gat;
  assign new_G378gat = ~G113gat | ~new_G290gat;
  assign new_G379gat = ~G120gat | ~new_G290gat;
  assign new_G380gat = ~G127gat | ~new_G293gat;
  assign new_G381gat = ~G134gat | ~new_G293gat;
  assign new_G382gat = ~G141gat | ~new_G296gat;
  assign new_G383gat = ~G148gat | ~new_G296gat;
  assign new_G384gat = ~G155gat | ~new_G299gat;
  assign new_G385gat = ~G162gat | ~new_G299gat;
  assign new_G386gat = ~G169gat | ~new_G302gat;
  assign new_G387gat = ~G176gat | ~new_G302gat;
  assign new_G388gat = ~G183gat | ~new_G305gat;
  assign new_G389gat = ~G190gat | ~new_G305gat;
  assign new_G390gat = ~G197gat | ~new_G308gat;
  assign new_G391gat = ~G204gat | ~new_G308gat;
  assign new_G392gat = ~G211gat | ~new_G311gat;
  assign new_G393gat = ~G218gat | ~new_G311gat;
  assign new_G394gat = ~G1gat | ~new_G314gat;
  assign new_G395gat = ~G29gat | ~new_G314gat;
  assign new_G396gat = ~G57gat | ~new_G317gat;
  assign new_G397gat = ~G85gat | ~new_G317gat;
  assign new_G398gat = ~G8gat | ~new_G320gat;
  assign new_G399gat = ~G36gat | ~new_G320gat;
  assign new_G400gat = ~G64gat | ~new_G323gat;
  assign new_G401gat = ~G92gat | ~new_G323gat;
  assign new_G402gat = ~G15gat | ~new_G326gat;
  assign new_G403gat = ~G43gat | ~new_G326gat;
  assign new_G404gat = ~G71gat | ~new_G329gat;
  assign new_G405gat = ~G99gat | ~new_G329gat;
  assign new_G406gat = ~G22gat | ~new_G332gat;
  assign new_G407gat = ~G50gat | ~new_G332gat;
  assign new_G408gat = ~G78gat | ~new_G335gat;
  assign new_G409gat = ~G106gat | ~new_G335gat;
  assign new_G410gat = ~G113gat | ~new_G338gat;
  assign new_G411gat = ~G141gat | ~new_G338gat;
  assign new_G412gat = ~G169gat | ~new_G341gat;
  assign new_G413gat = ~G197gat | ~new_G341gat;
  assign new_G414gat = ~G120gat | ~new_G344gat;
  assign new_G415gat = ~G148gat | ~new_G344gat;
  assign new_G416gat = ~G176gat | ~new_G347gat;
  assign new_G417gat = ~G204gat | ~new_G347gat;
  assign new_G418gat = ~G127gat | ~new_G350gat;
  assign new_G419gat = ~G155gat | ~new_G350gat;
  assign new_G420gat = ~G183gat | ~new_G353gat;
  assign new_G421gat = ~G211gat | ~new_G353gat;
  assign new_G422gat = ~G134gat | ~new_G356gat;
  assign new_G423gat = ~G162gat | ~new_G356gat;
  assign new_G424gat = ~G190gat | ~new_G359gat;
  assign new_G425gat = ~G218gat | ~new_G359gat;
  assign new_G426gat = ~new_G362gat | ~new_G363gat;
  assign new_G429gat = ~new_G364gat | ~new_G365gat;
  assign new_G432gat = ~new_G366gat | ~new_G367gat;
  assign new_G435gat = ~new_G368gat | ~new_G369gat;
  assign new_G438gat = ~new_G370gat | ~new_G371gat;
  assign new_G441gat = ~new_G372gat | ~new_G373gat;
  assign new_G444gat = ~new_G374gat | ~new_G375gat;
  assign new_G447gat = ~new_G376gat | ~new_G377gat;
  assign new_G450gat = ~new_G378gat | ~new_G379gat;
  assign new_G453gat = ~new_G380gat | ~new_G381gat;
  assign new_G456gat = ~new_G382gat | ~new_G383gat;
  assign new_G459gat = ~new_G384gat | ~new_G385gat;
  assign new_G462gat = ~new_G386gat | ~new_G387gat;
  assign new_G465gat = ~new_G388gat | ~new_G389gat;
  assign new_G468gat = ~new_G390gat | ~new_G391gat;
  assign new_G471gat = ~new_G392gat | ~new_G393gat;
  assign new_G474gat = ~new_G394gat | ~new_G395gat;
  assign new_G477gat = ~new_G396gat | ~new_G397gat;
  assign new_G480gat = ~new_G398gat | ~new_G399gat;
  assign new_G483gat = ~new_G400gat | ~new_G401gat;
  assign new_G486gat = ~new_G402gat | ~new_G403gat;
  assign new_G489gat = ~new_G404gat | ~new_G405gat;
  assign new_G492gat = ~new_G406gat | ~new_G407gat;
  assign new_G495gat = ~new_G408gat | ~new_G409gat;
  assign new_G498gat = ~new_G410gat | ~new_G411gat;
  assign new_G501gat = ~new_G412gat | ~new_G413gat;
  assign new_G504gat = ~new_G414gat | ~new_G415gat;
  assign new_G507gat = ~new_G416gat | ~new_G417gat;
  assign new_G510gat = ~new_G418gat | ~new_G419gat;
  assign new_G513gat = ~new_G420gat | ~new_G421gat;
  assign new_G516gat = ~new_G422gat | ~new_G423gat;
  assign new_G519gat = ~new_G424gat | ~new_G425gat;
  assign new_G522gat = ~new_G426gat | ~new_G429gat;
  assign new_G525gat = ~new_G432gat | ~new_G435gat;
  assign new_G528gat = ~new_G438gat | ~new_G441gat;
  assign new_G531gat = ~new_G444gat | ~new_G447gat;
  assign new_G534gat = ~new_G450gat | ~new_G453gat;
  assign new_G537gat = ~new_G456gat | ~new_G459gat;
  assign new_G540gat = ~new_G462gat | ~new_G465gat;
  assign new_G543gat = ~new_G468gat | ~new_G471gat;
  assign new_G546gat = ~new_G474gat | ~new_G477gat;
  assign new_G549gat = ~new_G480gat | ~new_G483gat;
  assign new_G552gat = ~new_G486gat | ~new_G489gat;
  assign new_G555gat = ~new_G492gat | ~new_G495gat;
  assign new_G558gat = ~new_G498gat | ~new_G501gat;
  assign new_G561gat = ~new_G504gat | ~new_G507gat;
  assign new_G564gat = ~new_G510gat | ~new_G513gat;
  assign new_G567gat = ~new_G516gat | ~new_G519gat;
  assign new_G570gat = ~new_G426gat | ~new_G522gat;
  assign new_G571gat = ~new_G429gat | ~new_G522gat;
  assign new_G572gat = ~new_G432gat | ~new_G525gat;
  assign new_G573gat = ~new_G435gat | ~new_G525gat;
  assign new_G574gat = ~new_G438gat | ~new_G528gat;
  assign new_G575gat = ~new_G441gat | ~new_G528gat;
  assign new_G576gat = ~new_G444gat | ~new_G531gat;
  assign new_G577gat = ~new_G447gat | ~new_G531gat;
  assign new_G578gat = ~new_G450gat | ~new_G534gat;
  assign new_G579gat = ~new_G453gat | ~new_G534gat;
  assign new_G580gat = ~new_G456gat | ~new_G537gat;
  assign new_G581gat = ~new_G459gat | ~new_G537gat;
  assign new_G582gat = ~new_G462gat | ~new_G540gat;
  assign new_G583gat = ~new_G465gat | ~new_G540gat;
  assign new_G584gat = ~new_G468gat | ~new_G543gat;
  assign new_G585gat = ~new_G471gat | ~new_G543gat;
  assign new_G586gat = ~new_G474gat | ~new_G546gat;
  assign new_G587gat = ~new_G477gat | ~new_G546gat;
  assign new_G588gat = ~new_G480gat | ~new_G549gat;
  assign new_G589gat = ~new_G483gat | ~new_G549gat;
  assign new_G590gat = ~new_G486gat | ~new_G552gat;
  assign new_G591gat = ~new_G489gat | ~new_G552gat;
  assign new_G592gat = ~new_G492gat | ~new_G555gat;
  assign new_G593gat = ~new_G495gat | ~new_G555gat;
  assign new_G594gat = ~new_G498gat | ~new_G558gat;
  assign new_G595gat = ~new_G501gat | ~new_G558gat;
  assign new_G596gat = ~new_G504gat | ~new_G561gat;
  assign new_G597gat = ~new_G507gat | ~new_G561gat;
  assign new_G598gat = ~new_G510gat | ~new_G564gat;
  assign new_G599gat = ~new_G513gat | ~new_G564gat;
  assign new_G600gat = ~new_G516gat | ~new_G567gat;
  assign new_G601gat = ~new_G519gat | ~new_G567gat;
  assign new_G602gat = ~new_G570gat | ~new_G571gat;
  assign new_G607gat = ~new_G572gat | ~new_G573gat;
  assign new_G612gat = ~new_G574gat | ~new_G575gat;
  assign new_G617gat = ~new_G576gat | ~new_G577gat;
  assign new_G622gat = ~new_G578gat | ~new_G579gat;
  assign new_G627gat = ~new_G580gat | ~new_G581gat;
  assign new_G632gat = ~new_G582gat | ~new_G583gat;
  assign new_G637gat = ~new_G584gat | ~new_G585gat;
  assign new_G642gat = ~new_G586gat | ~new_G587gat;
  assign new_G645gat = ~new_G588gat | ~new_G589gat;
  assign new_G648gat = ~new_G590gat | ~new_G591gat;
  assign new_G651gat = ~new_G592gat | ~new_G593gat;
  assign new_G654gat = ~new_G594gat | ~new_G595gat;
  assign new_G657gat = ~new_G596gat | ~new_G597gat;
  assign new_G660gat = ~new_G598gat | ~new_G599gat;
  assign new_G663gat = ~new_G600gat | ~new_G601gat;
  assign new_G666gat = ~new_G602gat | ~new_G607gat;
  assign new_G669gat = ~new_G612gat | ~new_G617gat;
  assign new_G672gat = ~new_G602gat | ~new_G612gat;
  assign new_G675gat = ~new_G607gat | ~new_G617gat;
  assign new_G678gat = ~new_G622gat | ~new_G627gat;
  assign new_G681gat = ~new_G632gat | ~new_G637gat;
  assign new_G684gat = ~new_G622gat | ~new_G632gat;
  assign new_G687gat = ~new_G627gat | ~new_G637gat;
  assign new_G690gat = ~new_G602gat | ~new_G666gat;
  assign new_G691gat = ~new_G607gat | ~new_G666gat;
  assign new_G692gat = ~new_G612gat | ~new_G669gat;
  assign new_G693gat = ~new_G617gat | ~new_G669gat;
  assign new_G694gat = ~new_G602gat | ~new_G672gat;
  assign new_G695gat = ~new_G612gat | ~new_G672gat;
  assign new_G696gat = ~new_G607gat | ~new_G675gat;
  assign new_G697gat = ~new_G617gat | ~new_G675gat;
  assign new_G698gat = ~new_G622gat | ~new_G678gat;
  assign new_G699gat = ~new_G627gat | ~new_G678gat;
  assign new_G700gat = ~new_G632gat | ~new_G681gat;
  assign new_G701gat = ~new_G637gat | ~new_G681gat;
  assign new_G702gat = ~new_G622gat | ~new_G684gat;
  assign new_G703gat = ~new_G632gat | ~new_G684gat;
  assign new_G704gat = ~new_G627gat | ~new_G687gat;
  assign new_G705gat = ~new_G637gat | ~new_G687gat;
  assign new_G706gat = ~new_G690gat | ~new_G691gat;
  assign new_G709gat = ~new_G692gat | ~new_G693gat;
  assign new_G712gat = ~new_G694gat | ~new_G695gat;
  assign new_G715gat = ~new_G696gat | ~new_G697gat;
  assign new_G718gat = ~new_G698gat | ~new_G699gat;
  assign new_G721gat = ~new_G700gat | ~new_G701gat;
  assign new_G724gat = ~new_G702gat | ~new_G703gat;
  assign new_G727gat = ~new_G704gat | ~new_G705gat;
  assign new_G730gat = ~new_G242gat | ~new_G718gat;
  assign new_G733gat = ~new_G245gat | ~new_G721gat;
  assign new_G736gat = ~new_G248gat | ~new_G724gat;
  assign new_G739gat = ~new_G251gat | ~new_G727gat;
  assign new_G742gat = ~new_G254gat | ~new_G706gat;
  assign new_G745gat = ~new_G257gat | ~new_G709gat;
  assign new_G748gat = ~new_G260gat | ~new_G712gat;
  assign new_G751gat = ~new_G263gat | ~new_G715gat;
  assign new_G754gat = ~new_G242gat | ~new_G730gat;
  assign new_G755gat = ~new_G718gat | ~new_G730gat;
  assign new_G756gat = ~new_G245gat | ~new_G733gat;
  assign new_G757gat = ~new_G721gat | ~new_G733gat;
  assign new_G758gat = ~new_G248gat | ~new_G736gat;
  assign new_G759gat = ~new_G724gat | ~new_G736gat;
  assign new_G760gat = ~new_G251gat | ~new_G739gat;
  assign new_G761gat = ~new_G727gat | ~new_G739gat;
  assign new_G762gat = ~new_G254gat | ~new_G742gat;
  assign new_G763gat = ~new_G706gat | ~new_G742gat;
  assign new_G764gat = ~new_G257gat | ~new_G745gat;
  assign new_G765gat = ~new_G709gat | ~new_G745gat;
  assign new_G766gat = ~new_G260gat | ~new_G748gat;
  assign new_G767gat = ~new_G712gat | ~new_G748gat;
  assign new_G768gat = ~new_G263gat | ~new_G751gat;
  assign new_G769gat = ~new_G715gat | ~new_G751gat;
  assign new_G770gat = ~new_G754gat | ~new_G755gat;
  assign new_G773gat = ~new_G756gat | ~new_G757gat;
  assign new_G776gat = ~new_G758gat | ~new_G759gat;
  assign new_G779gat = ~new_G760gat | ~new_G761gat;
  assign new_G782gat = ~new_G762gat | ~new_G763gat;
  assign new_G785gat = ~new_G764gat | ~new_G765gat;
  assign new_G788gat = ~new_G766gat | ~new_G767gat;
  assign new_G791gat = ~new_G768gat | ~new_G769gat;
  assign new_G794gat = ~new_G642gat | ~new_G770gat;
  assign new_G797gat = ~new_G645gat | ~new_G773gat;
  assign new_G800gat = ~new_G648gat | ~new_G776gat;
  assign new_G803gat = ~new_G651gat | ~new_G779gat;
  assign new_G806gat = ~new_G654gat | ~new_G782gat;
  assign new_G809gat = ~new_G657gat | ~new_G785gat;
  assign new_G812gat = ~new_G660gat | ~new_G788gat;
  assign new_G815gat = ~new_G663gat | ~new_G791gat;
  assign new_G818gat = ~new_G642gat | ~new_G794gat;
  assign new_G819gat = ~new_G770gat | ~new_G794gat;
  assign new_G820gat = ~new_G645gat | ~new_G797gat;
  assign new_G821gat = ~new_G773gat | ~new_G797gat;
  assign new_G822gat = ~new_G648gat | ~new_G800gat;
  assign new_G823gat = ~new_G776gat | ~new_G800gat;
  assign new_G824gat = ~new_G651gat | ~new_G803gat;
  assign new_G825gat = ~new_G779gat | ~new_G803gat;
  assign new_G826gat = ~new_G654gat | ~new_G806gat;
  assign new_G827gat = ~new_G782gat | ~new_G806gat;
  assign new_G828gat = ~new_G657gat | ~new_G809gat;
  assign new_G829gat = ~new_G785gat | ~new_G809gat;
  assign new_G830gat = ~new_G660gat | ~new_G812gat;
  assign new_G831gat = ~new_G788gat | ~new_G812gat;
  assign new_G832gat = ~new_G663gat | ~new_G815gat;
  assign new_G833gat = ~new_G791gat | ~new_G815gat;
  assign new_G834gat = ~new_G818gat | ~new_G819gat;
  assign new_G847gat = ~new_G820gat | ~new_G821gat;
  assign new_G860gat = ~new_G822gat | ~new_G823gat;
  assign new_G873gat = ~new_G824gat | ~new_G825gat;
  assign new_G886gat = ~new_G828gat | ~new_G829gat;
  assign new_G899gat = ~new_G832gat | ~new_G833gat;
  assign new_G912gat = ~new_G830gat | ~new_G831gat;
  assign new_G925gat = ~new_G826gat | ~new_G827gat;
  assign new_G938gat = ~new_G834gat;
  assign new_G939gat = ~new_G847gat;
  assign new_G940gat = ~new_G860gat;
  assign new_G941gat = ~new_G834gat;
  assign new_G942gat = ~new_G847gat;
  assign new_G943gat = ~new_G873gat;
  assign new_G944gat = ~new_G834gat;
  assign new_G945gat = ~new_G860gat;
  assign new_G946gat = ~new_G873gat;
  assign new_G947gat = ~new_G847gat;
  assign new_G948gat = ~new_G860gat;
  assign new_G949gat = ~new_G873gat;
  assign new_G950gat = ~new_G886gat;
  assign new_G951gat = ~new_G899gat;
  assign new_G952gat = ~new_G886gat;
  assign new_G953gat = ~new_G912gat;
  assign new_G954gat = ~new_G925gat;
  assign new_G955gat = ~new_G899gat;
  assign new_G956gat = ~new_G925gat;
  assign new_G957gat = ~new_G912gat;
  assign new_G958gat = ~new_G925gat;
  assign new_G959gat = ~new_G886gat;
  assign new_G960gat = ~new_G912gat;
  assign new_G961gat = ~new_G925gat;
  assign new_G962gat = ~new_G886gat;
  assign new_G963gat = ~new_G899gat;
  assign new_G964gat = ~new_G925gat;
  assign new_G965gat = ~new_G912gat;
  assign new_G966gat = ~new_G899gat;
  assign new_G967gat = ~new_G886gat;
  assign new_G968gat = ~new_G912gat;
  assign new_G969gat = ~new_G899gat;
  assign new_G970gat = ~new_G847gat;
  assign new_G971gat = ~new_G873gat;
  assign new_G972gat = ~new_G847gat;
  assign new_G973gat = ~new_G860gat;
  assign new_G974gat = ~new_G834gat;
  assign new_G975gat = ~new_G873gat;
  assign new_G976gat = ~new_G834gat;
  assign new_G977gat = ~new_G860gat;
  assign new_G978gat = new_G873gat & new_G940gat & new_G938gat & new_G939gat;
  assign new_G979gat = new_G943gat & new_G860gat & new_G941gat & new_G942gat;
  assign new_G980gat = new_G946gat & new_G945gat & new_G944gat & new_G847gat;
  assign new_G981gat = new_G949gat & new_G948gat & new_G834gat & new_G947gat;
  assign new_G982gat = new_G899gat & new_G960gat & new_G958gat & new_G959gat;
  assign new_G983gat = new_G963gat & new_G912gat & new_G961gat & new_G962gat;
  assign new_G984gat = new_G966gat & new_G965gat & new_G964gat & new_G886gat;
  assign new_G985gat = new_G969gat & new_G968gat & new_G925gat & new_G967gat;
  assign new_G986gat = new_G981gat | new_G980gat | new_G978gat | new_G979gat;
  assign new_G991gat = new_G985gat | new_G984gat | new_G982gat | new_G983gat;
  assign new_G996gat = new_G986gat & new_G951gat & new_G912gat & new_G925gat & new_G950gat;
  assign new_G1001gat = new_G986gat & new_G899gat & new_G953gat & new_G925gat & new_G952gat;
  assign new_G1006gat = new_G986gat & new_G955gat & new_G912gat & new_G954gat & new_G886gat;
  assign new_G1011gat = new_G986gat & new_G899gat & new_G957gat & new_G956gat & new_G886gat;
  assign new_G1016gat = new_G991gat & new_G971gat & new_G860gat & new_G834gat & new_G970gat;
  assign new_G1021gat = new_G991gat & new_G873gat & new_G973gat & new_G834gat & new_G972gat;
  assign new_G1026gat = new_G991gat & new_G975gat & new_G860gat & new_G974gat & new_G847gat;
  assign new_G1031gat = new_G991gat & new_G873gat & new_G977gat & new_G976gat & new_G847gat;
  assign new_G1036gat = new_G834gat & new_G996gat;
  assign new_G1039gat = new_G847gat & new_G996gat;
  assign new_G1042gat = new_G860gat & new_G996gat;
  assign new_G1045gat = new_G873gat & new_G996gat;
  assign new_G1048gat = new_G834gat & new_G1001gat;
  assign new_G1051gat = new_G847gat & new_G1001gat;
  assign new_G1054gat = new_G860gat & new_G1001gat;
  assign new_G1057gat = new_G873gat & new_G1001gat;
  assign new_G1060gat = new_G834gat & new_G1006gat;
  assign new_G1063gat = new_G847gat & new_G1006gat;
  assign new_G1066gat = new_G860gat & new_G1006gat;
  assign new_G1069gat = new_G873gat & new_G1006gat;
  assign new_G1072gat = new_G834gat & new_G1011gat;
  assign new_G1075gat = new_G847gat & new_G1011gat;
  assign new_G1078gat = new_G860gat & new_G1011gat;
  assign new_G1081gat = new_G873gat & new_G1011gat;
  assign new_G1084gat = new_G925gat & new_G1016gat;
  assign new_G1087gat = new_G886gat & new_G1016gat;
  assign new_G1090gat = new_G912gat & new_G1016gat;
  assign new_G1093gat = new_G899gat & new_G1016gat;
  assign new_G1096gat = new_G925gat & new_G1021gat;
  assign new_G1099gat = new_G886gat & new_G1021gat;
  assign new_G1102gat = new_G912gat & new_G1021gat;
  assign new_G1105gat = new_G899gat & new_G1021gat;
  assign new_G1108gat = new_G925gat & new_G1026gat;
  assign new_G1111gat = new_G886gat & new_G1026gat;
  assign new_G1114gat = new_G912gat & new_G1026gat;
  assign new_G1117gat = new_G899gat & new_G1026gat;
  assign new_G1120gat = new_G925gat & new_G1031gat;
  assign new_G1123gat = new_G886gat & new_G1031gat;
  assign new_G1126gat = new_G912gat & new_G1031gat;
  assign new_G1129gat = new_G899gat & new_G1031gat;
  assign new_G1132gat = ~G1gat | ~new_G1036gat;
  assign new_G1135gat = ~G8gat | ~new_G1039gat;
  assign new_G1138gat = ~G15gat | ~new_G1042gat;
  assign new_G1141gat = ~G22gat | ~new_G1045gat;
  assign new_G1144gat = ~G29gat | ~new_G1048gat;
  assign new_G1147gat = ~G36gat | ~new_G1051gat;
  assign new_G1150gat = ~G43gat | ~new_G1054gat;
  assign new_G1153gat = ~G50gat | ~new_G1057gat;
  assign new_G1156gat = ~G57gat | ~new_G1060gat;
  assign new_G1159gat = ~G64gat | ~new_G1063gat;
  assign new_G1162gat = ~G71gat | ~new_G1066gat;
  assign new_G1165gat = ~G78gat | ~new_G1069gat;
  assign new_G1168gat = ~G85gat | ~new_G1072gat;
  assign new_G1171gat = ~G92gat | ~new_G1075gat;
  assign new_G1174gat = ~G99gat | ~new_G1078gat;
  assign new_G1177gat = ~G106gat | ~new_G1081gat;
  assign new_G1180gat = ~G113gat | ~new_G1084gat;
  assign new_G1183gat = ~G120gat | ~new_G1087gat;
  assign new_G1186gat = ~G127gat | ~new_G1090gat;
  assign new_G1189gat = ~G134gat | ~new_G1093gat;
  assign new_G1192gat = ~G141gat | ~new_G1096gat;
  assign new_G1195gat = ~G148gat | ~new_G1099gat;
  assign new_G1198gat = ~G155gat | ~new_G1102gat;
  assign new_G1201gat = ~G162gat | ~new_G1105gat;
  assign new_G1204gat = ~G169gat | ~new_G1108gat;
  assign new_G1207gat = ~G176gat | ~new_G1111gat;
  assign new_G1210gat = ~G183gat | ~new_G1114gat;
  assign new_G1213gat = ~G190gat | ~new_G1117gat;
  assign new_G1216gat = ~G197gat | ~new_G1120gat;
  assign new_G1219gat = ~G204gat | ~new_G1123gat;
  assign new_G1222gat = ~G211gat | ~new_G1126gat;
  assign new_G1225gat = ~G218gat | ~new_G1129gat;
  assign new_G1228gat = ~G1gat | ~new_G1132gat;
  assign new_G1229gat = ~new_G1036gat | ~new_G1132gat;
  assign new_G1230gat = ~G8gat | ~new_G1135gat;
  assign new_G1231gat = ~new_G1039gat | ~new_G1135gat;
  assign new_G1232gat = ~G15gat | ~new_G1138gat;
  assign new_G1233gat = ~new_G1042gat | ~new_G1138gat;
  assign new_G1234gat = ~G22gat | ~new_G1141gat;
  assign new_G1235gat = ~new_G1045gat | ~new_G1141gat;
  assign new_G1236gat = ~G29gat | ~new_G1144gat;
  assign new_G1237gat = ~new_G1048gat | ~new_G1144gat;
  assign new_G1238gat = ~G36gat | ~new_G1147gat;
  assign new_G1239gat = ~new_G1051gat | ~new_G1147gat;
  assign new_G1240gat = ~G43gat | ~new_G1150gat;
  assign new_G1241gat = ~new_G1054gat | ~new_G1150gat;
  assign new_G1242gat = ~G50gat | ~new_G1153gat;
  assign new_G1243gat = ~new_G1057gat | ~new_G1153gat;
  assign new_G1244gat = ~G57gat | ~new_G1156gat;
  assign new_G1245gat = ~new_G1060gat | ~new_G1156gat;
  assign new_G1246gat = ~G64gat | ~new_G1159gat;
  assign new_G1247gat = ~new_G1063gat | ~new_G1159gat;
  assign new_G1248gat = ~G71gat | ~new_G1162gat;
  assign new_G1249gat = ~new_G1066gat | ~new_G1162gat;
  assign new_G1250gat = ~G78gat | ~new_G1165gat;
  assign new_G1251gat = ~new_G1069gat | ~new_G1165gat;
  assign new_G1252gat = ~G85gat | ~new_G1168gat;
  assign new_G1253gat = ~new_G1072gat | ~new_G1168gat;
  assign new_G1254gat = ~G92gat | ~new_G1171gat;
  assign new_G1255gat = ~new_G1075gat | ~new_G1171gat;
  assign new_G1256gat = ~G99gat | ~new_G1174gat;
  assign new_G1257gat = ~new_G1078gat | ~new_G1174gat;
  assign new_G1258gat = ~G106gat | ~new_G1177gat;
  assign new_G1259gat = ~new_G1081gat | ~new_G1177gat;
  assign new_G1260gat = ~G113gat | ~new_G1180gat;
  assign new_G1261gat = ~new_G1084gat | ~new_G1180gat;
  assign new_G1262gat = ~G120gat | ~new_G1183gat;
  assign new_G1263gat = ~new_G1087gat | ~new_G1183gat;
  assign new_G1264gat = ~G127gat | ~new_G1186gat;
  assign new_G1265gat = ~new_G1090gat | ~new_G1186gat;
  assign new_G1266gat = ~G134gat | ~new_G1189gat;
  assign new_G1267gat = ~new_G1093gat | ~new_G1189gat;
  assign new_G1268gat = ~G141gat | ~new_G1192gat;
  assign new_G1269gat = ~new_G1096gat | ~new_G1192gat;
  assign new_G1270gat = ~G148gat | ~new_G1195gat;
  assign new_G1271gat = ~new_G1099gat | ~new_G1195gat;
  assign new_G1272gat = ~G155gat | ~new_G1198gat;
  assign new_G1273gat = ~new_G1102gat | ~new_G1198gat;
  assign new_G1274gat = ~G162gat | ~new_G1201gat;
  assign new_G1275gat = ~new_G1105gat | ~new_G1201gat;
  assign new_G1276gat = ~G169gat | ~new_G1204gat;
  assign new_G1277gat = ~new_G1108gat | ~new_G1204gat;
  assign new_G1278gat = ~G176gat | ~new_G1207gat;
  assign new_G1279gat = ~new_G1111gat | ~new_G1207gat;
  assign new_G1280gat = ~G183gat | ~new_G1210gat;
  assign new_G1281gat = ~new_G1114gat | ~new_G1210gat;
  assign new_G1282gat = ~G190gat | ~new_G1213gat;
  assign new_G1283gat = ~new_G1117gat | ~new_G1213gat;
  assign new_G1284gat = ~G197gat | ~new_G1216gat;
  assign new_G1285gat = ~new_G1120gat | ~new_G1216gat;
  assign new_G1286gat = ~G204gat | ~new_G1219gat;
  assign new_G1287gat = ~new_G1123gat | ~new_G1219gat;
  assign new_G1288gat = ~G211gat | ~new_G1222gat;
  assign new_G1289gat = ~new_G1126gat | ~new_G1222gat;
  assign new_G1290gat = ~G218gat | ~new_G1225gat;
  assign new_G1291gat = ~new_G1129gat | ~new_G1225gat;
  assign new_G1292gat = ~new_G1228gat | ~new_G1229gat;
  assign new_G1293gat = ~new_G1230gat | ~new_G1231gat;
  assign new_G1294gat = ~new_G1232gat | ~new_G1233gat;
  assign new_G1295gat = ~new_G1234gat | ~new_G1235gat;
  assign new_G1296gat = ~new_G1236gat | ~new_G1237gat;
  assign new_G1297gat = ~new_G1238gat | ~new_G1239gat;
  assign new_G1298gat = ~new_G1240gat | ~new_G1241gat;
  assign new_G1299gat = ~new_G1242gat | ~new_G1243gat;
  assign new_G1300gat = ~new_G1244gat | ~new_G1245gat;
  assign new_G1301gat = ~new_G1246gat | ~new_G1247gat;
  assign new_G1302gat = ~new_G1248gat | ~new_G1249gat;
  assign new_G1303gat = ~new_G1250gat | ~new_G1251gat;
  assign new_G1304gat = ~new_G1252gat | ~new_G1253gat;
  assign new_G1305gat = ~new_G1254gat | ~new_G1255gat;
  assign new_G1306gat = ~new_G1256gat | ~new_G1257gat;
  assign new_G1307gat = ~new_G1258gat | ~new_G1259gat;
  assign new_G1308gat = ~new_G1260gat | ~new_G1261gat;
  assign new_G1309gat = ~new_G1262gat | ~new_G1263gat;
  assign new_G1310gat = ~new_G1264gat | ~new_G1265gat;
  assign new_G1311gat = ~new_G1266gat | ~new_G1267gat;
  assign new_G1312gat = ~new_G1268gat | ~new_G1269gat;
  assign new_G1313gat = ~new_G1270gat | ~new_G1271gat;
  assign new_G1314gat = ~new_G1272gat | ~new_G1273gat;
  assign new_G1315gat = ~new_G1274gat | ~new_G1275gat;
  assign new_G1316gat = ~new_G1276gat | ~new_G1277gat;
  assign new_G1317gat = ~new_G1278gat | ~new_G1279gat;
  assign new_G1318gat = ~new_G1280gat | ~new_G1281gat;
  assign new_G1319gat = ~new_G1282gat | ~new_G1283gat;
  assign new_G1320gat = ~new_G1284gat | ~new_G1285gat;
  assign new_G1321gat = ~new_G1286gat | ~new_G1287gat;
  assign new_G1322gat = ~new_G1288gat | ~new_G1289gat;
  assign new_G1323gat = ~new_G1290gat | ~new_G1291gat;
  assign G1324gat = new_G1292gat;
  assign G1325gat = new_G1293gat;
  assign G1326gat = new_G1294gat;
  assign G1327gat = new_G1295gat;
  assign G1328gat = new_G1296gat;
  assign G1329gat = new_G1297gat;
  assign G1330gat = new_G1298gat;
  assign G1331gat = new_G1299gat;
  assign G1332gat = new_G1300gat;
  assign G1333gat = new_G1301gat;
  assign G1334gat = new_G1302gat;
  assign G1335gat = new_G1303gat;
  assign G1336gat = new_G1304gat;
  assign G1337gat = new_G1305gat;
  assign G1338gat = new_G1306gat;
  assign G1339gat = new_G1307gat;
  assign G1340gat = new_G1308gat;
  assign G1341gat = new_G1309gat;
  assign G1342gat = new_G1310gat;
  assign G1343gat = new_G1311gat;
  assign G1344gat = new_G1312gat;
  assign G1345gat = new_G1313gat;
  assign G1346gat = new_G1314gat;
  assign G1347gat = new_G1315gat;
  assign G1348gat = new_G1316gat;
  assign G1349gat = new_G1317gat;
  assign G1350gat = new_G1318gat;
  assign G1351gat = new_G1319gat;
  assign G1352gat = new_G1320gat;
  assign G1353gat = new_G1321gat;
  assign G1354gat = new_G1322gat;
  assign G1355gat = new_G1323gat;
endmodule
