// Benchmark "./benchmarks/iscas85/c3540" written by ABC on Sun Apr 28 12:32:38 2024

module c3540  ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_G432, new_G442, new_G447, new_G456, new_G460, new_G463, new_G467,
    new_G476, new_G479, new_G483, new_G492, new_G501, new_G504, new_G513,
    new_G517, new_G526, new_G530, new_G540, new_G587, new_G704, new_G707,
    new_G714, new_G717, new_G724, new_G731, new_G732, new_G736, new_G741,
    new_G758, new_G776, new_G780, new_G788, new_G791, new_G798, new_G799,
    new_G802, new_G826, new_G828, new_G831, new_G833, new_G836, new_G839,
    new_G842, new_G845, new_G848, new_G851, new_G890, new_G898, new_G907,
    new_G1032, new_G1035, new_G1048, new_G1049, new_G1050, new_G1051,
    new_G1540, new_G1699, new_G1826, new_G1827, new_G1828, new_G2051,
    new_G2478, new_G2865, new_G2868, new_G2931, new_G2934, new_G2939,
    new_G2942, new_G2947, new_G2950, new_G2957, new_G2960, new_G3007,
    new_G3079, new_G3087, new_G3095, new_G3103, new_G3419, new_G588,
    new_G759, new_G1541, new_G1772, new_G1829, new_G1834, new_G2052,
    new_G625, new_G545, new_G546, new_G547, new_G548, new_G549, new_G550,
    new_G551, new_G552, new_G2937, new_G2938, new_G2945, new_G2946,
    new_G621, new_G626, new_G635, new_G636, new_G3085, new_G3101, new_G657,
    new_G675, new_G721, new_G784, new_G794, new_G807, new_G816, new_G823,
    new_G860, new_G861, new_G864, new_G893, new_G896, new_G897, new_G3093,
    new_G905, new_G906, new_G3109, new_G973, new_G980, new_G987, new_G994,
    new_G1001, new_G1008, new_G1015, new_G1022, new_G1038, new_G1043,
    new_G1054, new_G1057, new_G1512, new_G1681, new_G1717, new_G1724,
    new_G1731, new_G1738, new_G1745, new_G1752, new_G1759, new_G1766,
    new_G1773, new_G1790, new_G1808, new_G2278, new_G2481, new_G3425,
    new_G2871, new_G2874, new_G2953, new_G2954, new_G2963, new_G2964,
    new_G3010, new_G3013, new_G3017, new_G3020, new_G3027, new_G3030,
    new_G3037, new_G3040, new_G3082, new_G3090, new_G3098, new_G3106,
    new_G352, new_G553, new_G554, new_G555, new_G556, new_G560, new_G561,
    new_G650, new_G956, new_G974, new_G975, new_G976, new_G981, new_G982,
    new_G988, new_G989, new_G990, new_G995, new_G996, new_G997, new_G1002,
    new_G1003, new_G1004, new_G1009, new_G1010, new_G1016, new_G1017,
    new_G1018, new_G1023, new_G1024, new_G1025, new_G1720, new_G1727,
    new_G1734, new_G1741, new_G1748, new_G1755, new_G1762, new_G1769,
    new_G1791, new_G1809, new_G1851, new_G1901, new_G1952, new_G2002,
    new_G2057, new_G2109, new_G2162, new_G2214, new_G2955, new_G2956,
    new_G2965, new_G2966, new_G354, new_G557, new_G562, new_G586, new_G630,
    new_G634, new_G639, new_G642, new_G3086, new_G644, new_G646, new_G3102,
    new_G654, new_G660, new_G678, new_G804, new_G806, new_G855, new_G867,
    new_G903, new_G3094, new_G912, new_G3110, new_G915, new_G927, new_G941,
    new_G977, new_G978, new_G984, new_G985, new_G991, new_G992, new_G998,
    new_G999, new_G1005, new_G1006, new_G1012, new_G1013, new_G1019,
    new_G1020, new_G1026, new_G1027, new_G1060, new_G1063, new_G1066,
    new_G1069, new_G1527, new_G1530, new_G1542, new_G1563, new_G1572,
    new_G1581, new_G1585, new_G1589, new_G1593, new_G1597, new_G1601,
    new_G1605, new_G1716, new_G1718, new_G1723, new_G1725, new_G1730,
    new_G1732, new_G1737, new_G1739, new_G1744, new_G1746, new_G1751,
    new_G1753, new_G1758, new_G1760, new_G1765, new_G1767, new_G1852,
    new_G1856, new_G1870, new_G1902, new_G1906, new_G1920, new_G1953,
    new_G1957, new_G1971, new_G2003, new_G2007, new_G2021, new_G2058,
    new_G2062, new_G2076, new_G2110, new_G2114, new_G2128, new_G2163,
    new_G2167, new_G2181, new_G2215, new_G2219, new_G2233, new_G2285,
    new_G2288, new_G2289, new_G2293, new_G2298, new_G2302, new_G2877,
    new_G2983, new_G2986, new_G3014, new_G3015, new_G3023, new_G3024,
    new_G3033, new_G3034, new_G3043, new_G3044, new_G643, new_G647,
    new_G680, new_G904, new_G913, new_G920, new_G979, new_G993, new_G1000,
    new_G1007, new_G1021, new_G1028, new_G1719, new_G1721, new_G1726,
    new_G1728, new_G1733, new_G1735, new_G1740, new_G1742, new_G1747,
    new_G1749, new_G1754, new_G1756, new_G1761, new_G1763, new_G1768,
    new_G1770, new_G1794, new_G1799, new_G1812, new_G1817, new_G1859,
    new_G1909, new_G1960, new_G2010, new_G2065, new_G2117, new_G2170,
    new_G2222, new_G2678, new_G2697, new_G2716, new_G2733, new_G2751,
    new_G2768, new_G2785, new_G2802, new_G3016, new_G3025, new_G3026,
    new_G3035, new_G3036, new_G3045, new_G3046, new_G2989, new_G2990,
    new_G610, new_G613, new_G616, new_G640, new_G648, new_G655, new_G665,
    new_G668, new_G671, new_G683, new_G685, new_G688, new_G694, new_G696,
    new_G699, new_G870, new_G887, new_G901, new_G910, new_G914, new_G916,
    new_G942, new_G943, new_G1072, new_G1084, new_G1096, new_G1108,
    new_G1120, new_G1132, new_G1144, new_G1156, new_G1533, new_G1534,
    new_G1535, new_G1545, new_G1554, new_G1610, new_G1619, new_G1628,
    new_G1637, new_G1646, new_G1655, new_G1664, new_G1673, new_G1722,
    new_G1729, new_G1736, new_G1743, new_G1750, new_G1757, new_G1764,
    new_G1771, new_G1853, new_G1954, new_G2004, new_G2059, new_G2164,
    new_G2216, new_G2485, new_G2900, new_G2903, new_G2967, new_G2970,
    new_G2975, new_G2978, new_G3047, new_G3050, new_G3055, new_G3058,
    new_G574, new_G575, new_G617, new_G641, new_G649, new_G662, new_G672,
    new_G690, new_G691, new_G701, new_G702, new_G902, new_G911, new_G917,
    new_G923, new_G1538, new_G1871, new_G1872, new_G1873, new_G1921,
    new_G1922, new_G1923, new_G1972, new_G1973, new_G1974, new_G2022,
    new_G2023, new_G2024, new_G2077, new_G2078, new_G2079, new_G2129,
    new_G2130, new_G2131, new_G2182, new_G2183, new_G2184, new_G2234,
    new_G2235, new_G2236, new_G2973, new_G2974, new_G2981, new_G2982,
    new_G576, new_G3053, new_G3054, new_G3061, new_G3062, new_G645,
    new_G926, new_G928, new_G947, new_G983, new_G1011, new_G1075,
    new_G1087, new_G1099, new_G1111, new_G1123, new_G1135, new_G1147,
    new_G1159, new_G1168, new_G1177, new_G1186, new_G1195, new_G1204,
    new_G1213, new_G1222, new_G1231, new_G1609, new_G1611, new_G1618,
    new_G1620, new_G1627, new_G1629, new_G1636, new_G1638, new_G1645,
    new_G1647, new_G1654, new_G1656, new_G1663, new_G1665, new_G1672,
    new_G1674, new_G1862, new_G1866, new_G1874, new_G1924, new_G1963,
    new_G1967, new_G1975, new_G2013, new_G2017, new_G2025, new_G2068,
    new_G2072, new_G2080, new_G2132, new_G2173, new_G2177, new_G2185,
    new_G2225, new_G2229, new_G2237, new_G2488, new_G2679, new_G2680,
    new_G2698, new_G2699, new_G2717, new_G2718, new_G2734, new_G2735,
    new_G2752, new_G2753, new_G2769, new_G2770, new_G2786, new_G2787,
    new_G2803, new_G2804, new_G359, new_G1029, new_G565, new_G566,
    new_G569, new_G570, new_G589, new_G590, new_G595, new_G596, new_G929,
    new_G938, new_G944, new_G986, new_G1014, new_G1616, new_G1625,
    new_G1634, new_G1643, new_G360, new_G567, new_G571, new_G579, new_G591,
    new_G597, new_G614, new_G1240, new_G1241, new_G1242, new_G1243,
    new_G1244, new_G1245, new_G1246, new_G1247, new_G1257, new_G1258,
    new_G1259, new_G1260, new_G1261, new_G1262, new_G1263, new_G1264,
    new_G1274, new_G1275, new_G1276, new_G1277, new_G1278, new_G1279,
    new_G1280, new_G1281, new_G1291, new_G1292, new_G1293, new_G1294,
    new_G1295, new_G1296, new_G1297, new_G1298, new_G1308, new_G1309,
    new_G1310, new_G1311, new_G1312, new_G1313, new_G1314, new_G1315,
    new_G1325, new_G1326, new_G1327, new_G1328, new_G1329, new_G1330,
    new_G1331, new_G1332, new_G1342, new_G1343, new_G1344, new_G1345,
    new_G1346, new_G1347, new_G1348, new_G1349, new_G1359, new_G1360,
    new_G1361, new_G1362, new_G1363, new_G1364, new_G1365, new_G1366,
    new_G1376, new_G1377, new_G1378, new_G1379, new_G1380, new_G1381,
    new_G1382, new_G1383, new_G1393, new_G1394, new_G1395, new_G1396,
    new_G1397, new_G1398, new_G1399, new_G1400, new_G1410, new_G1411,
    new_G1412, new_G1413, new_G1414, new_G1415, new_G1416, new_G1417,
    new_G1427, new_G1428, new_G1429, new_G1430, new_G1431, new_G1432,
    new_G1433, new_G1434, new_G1444, new_G1445, new_G1446, new_G1447,
    new_G1448, new_G1449, new_G1450, new_G1451, new_G1461, new_G1462,
    new_G1463, new_G1464, new_G1465, new_G1466, new_G1467, new_G1468,
    new_G1478, new_G1479, new_G1480, new_G1481, new_G1482, new_G1483,
    new_G1484, new_G1485, new_G1495, new_G1496, new_G1497, new_G1498,
    new_G1499, new_G1500, new_G1501, new_G1502, new_G1877, new_G1880,
    new_G1891, new_G1903, new_G1927, new_G1930, new_G1978, new_G1981,
    new_G1992, new_G2028, new_G2031, new_G2042, new_G2085, new_G2088,
    new_G2099, new_G2111, new_G2137, new_G2140, new_G2190, new_G2193,
    new_G2204, new_G2242, new_G2245, new_G2256, new_G2320, new_G2341,
    new_G2354, new_G2367, new_G2383, new_G2391, new_G2474, new_G2475,
    new_G2476, new_G2477, new_G2482, new_G568, new_G618, new_G1248,
    new_G1249, new_G1250, new_G1251, new_G1252, new_G1253, new_G1254,
    new_G1255, new_G1265, new_G1266, new_G1267, new_G1268, new_G1269,
    new_G1270, new_G1271, new_G1272, new_G1282, new_G1283, new_G1284,
    new_G1285, new_G1286, new_G1287, new_G1288, new_G1289, new_G1299,
    new_G1300, new_G1301, new_G1302, new_G1303, new_G1304, new_G1305,
    new_G1306, new_G1316, new_G1317, new_G1318, new_G1319, new_G1320,
    new_G1321, new_G1322, new_G1323, new_G1333, new_G1334, new_G1335,
    new_G1336, new_G1337, new_G1338, new_G1339, new_G1340, new_G1350,
    new_G1351, new_G1352, new_G1353, new_G1354, new_G1355, new_G1356,
    new_G1357, new_G1367, new_G1368, new_G1369, new_G1370, new_G1371,
    new_G1372, new_G1373, new_G1374, new_G1384, new_G1385, new_G1386,
    new_G1387, new_G1388, new_G1389, new_G1390, new_G1391, new_G1401,
    new_G1402, new_G1403, new_G1404, new_G1405, new_G1406, new_G1407,
    new_G1408, new_G1418, new_G1419, new_G1420, new_G1421, new_G1422,
    new_G1423, new_G1424, new_G1425, new_G1435, new_G1436, new_G1437,
    new_G1438, new_G1439, new_G1440, new_G1441, new_G1442, new_G1452,
    new_G1453, new_G1454, new_G1455, new_G1456, new_G1457, new_G1458,
    new_G1459, new_G1469, new_G1470, new_G1471, new_G1472, new_G1473,
    new_G1474, new_G1475, new_G1476, new_G1486, new_G1487, new_G1488,
    new_G1489, new_G1490, new_G1491, new_G1492, new_G1493, new_G1503,
    new_G1504, new_G1505, new_G1506, new_G1507, new_G1508, new_G1509,
    new_G1510, new_G2483, new_G600, new_G661, new_G669, new_G679,
    new_G1256, new_G1273, new_G1290, new_G1307, new_G1324, new_G1341,
    new_G1358, new_G1375, new_G1392, new_G1409, new_G1426, new_G1443,
    new_G1460, new_G1477, new_G1494, new_G1511, new_G1652, new_G1883,
    new_G1886, new_G1889, new_G1890, new_G1912, new_G1916, new_G1984,
    new_G1987, new_G1990, new_G1991, new_G2034, new_G2037, new_G2040,
    new_G2041, new_G2091, new_G2094, new_G2097, new_G2098, new_G2120,
    new_G2124, new_G2196, new_G2199, new_G2202, new_G2203, new_G2248,
    new_G2251, new_G2254, new_G2255, new_G2484, new_G2991, new_G2994,
    new_G2999, new_G3002, new_G3063, new_G3071, new_G3124, new_G3134,
    new_G3158, new_G3166, new_G3174, new_G3182, new_G3190, new_G3200,
    new_G3224, new_G3232, new_G3240, new_G3248, new_G663, new_G673,
    new_G681, new_G1536, new_G1537, new_G1582, new_G1583, new_G1586,
    new_G1587, new_G1590, new_G1591, new_G1594, new_G1595, new_G1598,
    new_G1599, new_G1602, new_G1603, new_G1606, new_G1607, new_G1894,
    new_G1997, new_G2047, new_G2102, new_G2209, new_G2261, new_G2489,
    new_G3005, new_G3006, new_G3077, new_G3069, new_G2997, new_G2998,
    new_G689, new_G700, new_G1539, new_G1584, new_G1588, new_G1592,
    new_G1596, new_G1600, new_G1604, new_G1608, new_G1661, new_G1892,
    new_G1893, new_G1933, new_G1936, new_G1939, new_G1940, new_G1941,
    new_G1993, new_G1996, new_G2043, new_G2046, new_G2100, new_G2101,
    new_G2143, new_G2146, new_G2149, new_G2150, new_G2151, new_G2205,
    new_G2208, new_G2257, new_G2260, new_G3138, new_G2328, new_G3162,
    new_G3170, new_G3178, new_G3186, new_G3204, new_G2375, new_G3236,
    new_G3244, new_G3252, new_G3228, new_G3066, new_G3074, new_G3128,
    new_G3194, new_G619, new_G620, new_G582, new_G583, new_G692, new_G703,
    new_G1612, new_G1621, new_G1630, new_G1639, new_G1648, new_G1657,
    new_G1666, new_G1675, new_G1895, new_G1946, new_G1998, new_G2048,
    new_G2103, new_G2156, new_G2210, new_G2262, new_G2271, new_G2311,
    new_G356, new_G357, new_G603, new_G3078, new_G606, new_G3070,
    new_G1670, new_G1679, new_G1942, new_G1945, new_G2152, new_G2155,
    new_G2445, new_G2448, new_G2455, new_G2458, new_G3142, new_G3150,
    new_G3208, new_G3216, new_G604, new_G607, new_G1947, new_G2157,
    new_G2317, new_G2338, new_G2351, new_G2364, new_G2380, new_G2388,
    new_G605, new_G608, new_G2272, new_G2312, new_G3146, new_G3154,
    new_G3220, new_G3212, new_G2444, new_G2451, new_G2454, new_G2461,
    new_G2530, new_G3323, new_G349, new_G350, new_G2265, new_G2273,
    new_G2274, new_G2309, new_G2313, new_G2314, new_G2325, new_G2372,
    new_G2523, new_G2533, new_G3121, new_G3131, new_G3155, new_G3163,
    new_G3171, new_G3179, new_G3187, new_G3197, new_G3221, new_G3229,
    new_G3237, new_G3245, new_G2275, new_G2315, new_G3329, new_G2324,
    new_G2350, new_G2363, new_G2371, new_G2387, new_G2400, new_G2268,
    new_G3137, new_G3161, new_G2345, new_G3169, new_G3177, new_G2358,
    new_G3185, new_G3203, new_G3235, new_G3243, new_G2395, new_G3251,
    new_G3227, new_G2432, new_G2490, new_G3127, new_G3130, new_G3139,
    new_G3147, new_G3193, new_G3196, new_G3205, new_G3213, new_G2307,
    new_G2308, new_G2323, new_G2349, new_G2362, new_G2370, new_G2386,
    new_G2399, new_G2344, new_G2357, new_G2394, new_G2431, new_G2464,
    new_G2491, new_G3129, new_G3195, new_G368, new_G1615, new_G2337,
    new_G1633, new_G1642, new_G1651, new_G2379, new_G1669, new_G1678,
    new_G3145, new_G2332, new_G3153, new_G2346, new_G2359, new_G3219,
    new_G2396, new_G3211, new_G2425, new_G2433, new_G3272, new_G3308,
    new_G1613, new_G2336, new_G1631, new_G1640, new_G1649, new_G2378,
    new_G1667, new_G1676, new_G2331, new_G2424, new_G2467, new_G2495,
    new_G3295, new_G3374, new_G1614, new_G1624, new_G1632, new_G1641,
    new_G1650, new_G1660, new_G1668, new_G1677, new_G2333, new_G2406,
    new_G2409, new_G2415, new_G2419, new_G2426, new_G2439, new_G2518,
    new_G3276, new_G3312, new_G2612, new_G3326, new_G1617, new_G1622,
    new_G1635, new_G1644, new_G1653, new_G1658, new_G1671, new_G1680,
    new_G2500, new_G2505, new_G2519, new_G3378, new_G2642, new_G2645,
    new_G3301, new_G1623, new_G1659, new_G2401, new_G2501, new_G2511,
    new_G2512, new_G2513, new_G2514, new_G2517, new_G2531, new_G2532,
    new_G2534, new_G2535, new_G2607, new_G3330, new_G2643, new_G2687,
    new_G2725, new_G2742, new_G2760, new_G2794, new_G2811, new_G3280,
    new_G3290, new_G3298, new_G3316, new_G3406, new_G3414, new_G3422,
    new_G1626, new_G1662, new_G2567, new_G2589, new_G2608, new_G2654,
    new_G3253, new_G3277, new_G3287, new_G3305, new_G3313, new_G3350,
    new_G932, new_G2508, new_G2524, new_G2525, new_G2526, new_G3294,
    new_G2609, new_G3410, new_G3418, new_G2624, new_G3426, new_G2629,
    new_G2647, new_G2706, new_G2777, new_G3264, new_G3284, new_G3302,
    new_G3303, new_G3320, new_G3398, new_G2657, new_G398, new_G933,
    new_G2527, new_G3259, new_G3354, new_G3293, new_G2563, new_G3311,
    new_G2585, new_G2625, new_G3283, new_G3286, new_G3304, new_G3319,
    new_G3322, new_G3358, new_G3366, new_G3382, new_G3390, new_G397,
    new_G2544, new_G2562, new_G2584, new_G3402, new_G2626, new_G2632,
    new_G2634, new_G2650, new_G3268, new_G3256, new_G3285, new_G3321,
    new_G3371, new_G3403, new_G3411, new_G362, new_G1030, new_G2564,
    new_G3362, new_G3370, new_G2586, new_G3386, new_G3394, new_G2633,
    new_G3261, new_G3269, new_G3347, new_G3395, new_G363, new_G2536,
    new_G3260, new_G3377, new_G2580, new_G3409, new_G2616, new_G3417,
    new_G2622, new_G2635, new_G2805, new_G2808, new_G3334, new_G3342,
    new_G3454, new_G2537, new_G3275, new_G2540, new_G3353, new_G2557,
    new_G2579, new_G3401, new_G2602, new_G2615, new_G2621, new_G3267,
    new_G3112, new_G3355, new_G3363, new_G3379, new_G3387, new_G2538,
    new_G2539, new_G3338, new_G3346, new_G2556, new_G2581, new_G2601,
    new_G2617, new_G2623, new_G2638, new_G3458, new_G2814, new_G2816,
    new_G3111, new_G2541, new_G2558, new_G3361, new_G2571, new_G3369,
    new_G2577, new_G3385, new_G2593, new_G3393, new_G2598, new_G2603,
    new_G3113, new_G3116, new_G3451, new_G395, new_G2570, new_G2576,
    new_G2592, new_G2597, new_G2736, new_G2739, new_G2788, new_G3438,
    new_G3446, new_G3459, new_G3119, new_G3120, new_G2572, new_G2578,
    new_G2594, new_G2599, new_G2677, new_G3457, new_G2700, new_G2771,
    new_G3331, new_G3339, new_G3427, new_G3443, new_G954, new_G955,
    new_G2600, new_G3442, new_G3450, new_G2676, new_G2745, new_G2748,
    new_G3465, new_G3435, new_G950, new_G3337, new_G2548, new_G3345,
    new_G2553, new_G2661, new_G2662, new_G3433, new_G3449, new_G2672,
    new_G2674, new_G2719, new_G2754, new_G3430, new_G383, new_G951,
    new_G2547, new_G2552, new_G2663, new_G2670, new_G3441, new_G2671,
    new_G2675, new_G3491, new_G3499, new_G2549, new_G2554, new_G2664,
    new_G3434, new_G2669, new_G2673, new_G2757, new_G2791, new_G365,
    new_G1031, new_G2555, new_G2665, new_G2667, new_G2774, new_G3497,
    new_G3505, new_G366, new_G2658, new_G2659, new_G2666, new_G2668,
    new_G2681, new_G2763, new_G2765, new_G2797, new_G2799, new_G2660,
    new_G2703, new_G2722, new_G2780, new_G2782, new_G386, new_G392,
    new_G2684, new_G3462, new_G3470, new_G389, new_G2709, new_G2713,
    new_G2728, new_G2730, new_G2922, new_G3467, new_G2690, new_G2694,
    new_G2821, new_G3466, new_G3474, new_G380, new_G2822, new_G3473,
    new_G2827, new_G2839, new_G2883, new_G3507, new_G2823, new_G2826,
    new_G2880, new_G2925, new_G2928, new_G3510, new_G2828, new_G3494,
    new_G3502, new_G3513, new_G3544, new_G3552, new_G406, new_G2929,
    new_G3475, new_G3483, new_G3514, new_G3515, new_G3541, new_G3549,
    new_G2930, new_G2842, new_G3498, new_G2852, new_G3506, new_G3548,
    new_G3556, new_G3478, new_G3486, new_G3516, new_G408, new_G3481,
    new_G3489, new_G2843, new_G2853, new_G3547, new_G2887, new_G2896,
    new_G3555, new_G3520, new_G2831, new_G3482, new_G2836, new_G3490,
    new_G2844, new_G2848, new_G2886, new_G2895, new_G2832, new_G2837,
    new_G2849, new_G3524, new_G2888, new_G2891, new_G2833, new_G2838,
    new_G2892, new_G3517, new_G2906, new_G2908, new_G2913, new_G3523,
    new_G2855, new_G2907, new_G2909, new_G3525, new_G3533, new_G2854,
    new_G2910, new_G3560, new_G3568, new_G2856, new_G3539, new_G3531,
    new_G3572, new_G3564, new_G3557, new_G3565, new_G3528, new_G3536,
    new_G2921, new_G2917, new_G3571, new_G3563, new_G2863, new_G2859,
    new_G2920, new_G2916, new_G3540, new_G3532, new_G2864, new_G2860,
    new_G403, new_G404, new_G400, new_G401;
  assign new_G432 = G50;
  assign new_G442 = ~G50;
  assign new_G447 = G58;
  assign new_G456 = ~G58;
  assign new_G460 = G68;
  assign new_G463 = ~G68;
  assign new_G467 = G68;
  assign new_G476 = G77;
  assign new_G479 = ~G77;
  assign new_G483 = G77;
  assign new_G492 = G87;
  assign new_G501 = ~G87;
  assign new_G504 = G97;
  assign new_G513 = ~G97;
  assign new_G517 = G107;
  assign new_G526 = ~G107;
  assign new_G530 = G116;
  assign new_G540 = ~G116;
  assign new_G587 = G257 | G264;
  assign new_G704 = ~G1;
  assign new_G707 = G1;
  assign new_G714 = ~G1;
  assign new_G717 = G13;
  assign new_G724 = ~G13;
  assign new_G731 = G13 & G20;
  assign new_G732 = ~G20;
  assign new_G736 = G20;
  assign new_G741 = ~G20;
  assign new_G758 = ~G33;
  assign new_G776 = G33;
  assign new_G780 = ~G33;
  assign new_G788 = G33 & G41;
  assign new_G791 = ~G41;
  assign new_G798 = G41 | G45;
  assign new_G799 = G45;
  assign new_G802 = ~G45;
  assign new_G826 = ~G50;
  assign new_G828 = G58;
  assign new_G831 = ~G58;
  assign new_G833 = G68;
  assign new_G836 = ~G68;
  assign new_G839 = G87;
  assign new_G842 = ~G87;
  assign new_G845 = G97;
  assign new_G848 = ~G97;
  assign new_G851 = ~G107;
  assign new_G890 = G1;
  assign new_G898 = G68;
  assign new_G907 = G107;
  assign new_G1032 = ~G20;
  assign new_G1035 = G190;
  assign new_G1048 = ~G200;
  assign new_G1049 = G20 & G200;
  assign new_G1050 = ~G20 | ~G200;
  assign new_G1051 = G20 & G179;
  assign new_G1540 = ~G20;
  assign new_G1699 = G1698 | G33;
  assign new_G1826 = ~G1 | ~G13;
  assign new_G1827 = ~G33 | ~G1 | ~G20;
  assign new_G1828 = ~G20;
  assign new_G2051 = ~G33;
  assign new_G2478 = G179;
  assign new_G2865 = ~G213;
  assign new_G2868 = G343;
  assign new_G2931 = G226;
  assign new_G2934 = G232;
  assign new_G2939 = G238;
  assign new_G2942 = G244;
  assign new_G2947 = G250;
  assign new_G2950 = G257;
  assign new_G2957 = G264;
  assign new_G2960 = G270;
  assign new_G3007 = G50;
  assign new_G3079 = G58;
  assign new_G3087 = G58;
  assign new_G3095 = G97;
  assign new_G3103 = G97;
  assign new_G3419 = G330;
  assign new_G588 = G250 & new_G587;
  assign new_G759 = new_G758 | G20;
  assign new_G1541 = new_G1540 | G169;
  assign new_G1772 = ~new_G731;
  assign new_G1829 = new_G1828 | G1;
  assign new_G1834 = new_G1826 & new_G1827;
  assign new_G2052 = new_G2051 | G1;
  assign new_G625 = new_G836 & new_G826 & new_G831;
  assign new_G545 = ~G226 | ~new_G432;
  assign new_G546 = ~G232 | ~new_G447;
  assign new_G547 = ~G238 | ~new_G467;
  assign new_G548 = ~G244 | ~new_G483;
  assign new_G549 = ~G250 | ~new_G492;
  assign new_G550 = ~G257 | ~new_G504;
  assign new_G551 = ~G264 | ~new_G517;
  assign new_G552 = ~G270 | ~new_G530;
  assign new_G2937 = ~new_G2931;
  assign new_G2938 = ~new_G2934;
  assign new_G2945 = ~new_G2939;
  assign new_G2946 = ~new_G2942;
  assign new_G621 = ~new_G456 | ~new_G463;
  assign new_G626 = ~new_G513 | ~new_G526;
  assign new_G635 = ~new_G460 | ~new_G476;
  assign new_G636 = new_G442;
  assign new_G3085 = ~new_G3079;
  assign new_G3101 = ~new_G3095;
  assign new_G657 = new_G802;
  assign new_G675 = new_G802;
  assign new_G721 = new_G717;
  assign new_G784 = new_G780;
  assign new_G794 = new_G791;
  assign new_G807 = new_G714 & new_G798;
  assign new_G816 = new_G791 & new_G714 & new_G799;
  assign new_G823 = new_G704 & new_G799;
  assign new_G860 = new_G736 & new_G707 & new_G724;
  assign new_G861 = ~new_G736 | ~new_G707 | ~new_G724;
  assign new_G864 = ~new_G707 | ~new_G724;
  assign new_G893 = new_G890;
  assign new_G896 = ~G45 | ~new_G717 | ~new_G732;
  assign new_G897 = ~new_G836 | ~new_G826 | ~new_G831;
  assign new_G3093 = ~new_G3087;
  assign new_G905 = new_G851 & new_G842 & new_G848;
  assign new_G906 = ~new_G851 | ~new_G842 | ~new_G848;
  assign new_G3109 = ~new_G3103;
  assign new_G973 = ~new_G741;
  assign new_G980 = ~new_G741;
  assign new_G987 = ~new_G741;
  assign new_G994 = ~new_G741;
  assign new_G1001 = ~new_G741;
  assign new_G1008 = ~new_G741;
  assign new_G1015 = ~new_G741;
  assign new_G1022 = ~new_G741;
  assign new_G1038 = new_G1032 | new_G1035;
  assign new_G1043 = ~new_G1032 & ~new_G1035;
  assign new_G1054 = new_G1051;
  assign new_G1057 = ~new_G1051;
  assign new_G1512 = new_G776;
  assign new_G1681 = new_G780;
  assign new_G1717 = ~new_G1699;
  assign new_G1724 = ~new_G1699;
  assign new_G1731 = ~new_G1699;
  assign new_G1738 = ~new_G1699;
  assign new_G1745 = ~new_G1699;
  assign new_G1752 = ~new_G1699;
  assign new_G1759 = ~new_G1699;
  assign new_G1766 = ~new_G1699;
  assign new_G1773 = G1 | new_G1772;
  assign new_G1790 = ~new_G788;
  assign new_G1808 = ~new_G788;
  assign new_G2278 = new_G732 & new_G704 & new_G717;
  assign new_G2481 = ~new_G2478;
  assign new_G3425 = ~new_G3419;
  assign new_G2871 = new_G2865 | new_G2868;
  assign new_G2874 = ~new_G2865 & ~new_G2868;
  assign new_G2953 = ~new_G2947;
  assign new_G2954 = ~new_G2950;
  assign new_G2963 = ~new_G2957;
  assign new_G2964 = ~new_G2960;
  assign new_G3010 = new_G456;
  assign new_G3013 = ~new_G3007;
  assign new_G3017 = new_G463;
  assign new_G3020 = new_G479;
  assign new_G3027 = new_G501;
  assign new_G3030 = new_G513;
  assign new_G3037 = new_G526;
  assign new_G3040 = new_G540;
  assign new_G3082 = new_G898;
  assign new_G3090 = new_G898;
  assign new_G3098 = new_G907;
  assign new_G3106 = new_G907;
  assign new_G352 = ~new_G479 | ~new_G625;
  assign new_G553 = new_G548 & new_G547 & new_G545 & new_G546;
  assign new_G554 = new_G552 & new_G551 & new_G549 & new_G550;
  assign new_G555 = ~new_G2934 | ~new_G2937;
  assign new_G556 = ~new_G2931 | ~new_G2938;
  assign new_G560 = ~new_G2942 | ~new_G2945;
  assign new_G561 = ~new_G2939 | ~new_G2946;
  assign new_G650 = new_G432 & new_G621;
  assign new_G956 = new_G890 & new_G896;
  assign new_G974 = ~new_G759;
  assign new_G975 = new_G741 & new_G759;
  assign new_G976 = new_G897 & new_G973;
  assign new_G981 = ~new_G759;
  assign new_G982 = new_G741 & new_G759;
  assign new_G988 = ~new_G759;
  assign new_G989 = new_G741 & new_G759;
  assign new_G990 = new_G836 & new_G987;
  assign new_G995 = ~new_G759;
  assign new_G996 = new_G741 & new_G759;
  assign new_G997 = G77 & new_G994;
  assign new_G1002 = ~new_G759;
  assign new_G1003 = new_G741 & new_G759;
  assign new_G1004 = new_G906 & new_G1001;
  assign new_G1009 = ~new_G759;
  assign new_G1010 = new_G741 & new_G759;
  assign new_G1016 = ~new_G759;
  assign new_G1017 = new_G741 & new_G759;
  assign new_G1018 = new_G851 & new_G1015;
  assign new_G1023 = ~new_G759;
  assign new_G1024 = new_G741 & new_G759;
  assign new_G1025 = G116 & new_G1022;
  assign new_G1720 = G222 & new_G1717;
  assign new_G1727 = G223 & new_G1724;
  assign new_G1734 = G226 & new_G1731;
  assign new_G1741 = G232 & new_G1738;
  assign new_G1748 = G238 & new_G1745;
  assign new_G1755 = G244 & new_G1752;
  assign new_G1762 = G250 & new_G1759;
  assign new_G1769 = G257 & new_G1766;
  assign new_G1791 = new_G1790 & G1 & G13;
  assign new_G1809 = new_G1808 & G1 & G13;
  assign new_G1851 = ~new_G1834;
  assign new_G1901 = ~new_G1834;
  assign new_G1952 = ~new_G1834;
  assign new_G2002 = ~new_G1834;
  assign new_G2057 = ~new_G1834;
  assign new_G2109 = ~new_G1834;
  assign new_G2162 = ~new_G1834;
  assign new_G2214 = ~new_G1834;
  assign new_G2955 = ~new_G2950 | ~new_G2953;
  assign new_G2956 = ~new_G2947 | ~new_G2954;
  assign new_G2965 = ~new_G2960 | ~new_G2963;
  assign new_G2966 = ~new_G2957 | ~new_G2964;
  assign G353 = ~new_G352;
  assign new_G354 = G87 & new_G626;
  assign new_G557 = ~new_G555 | ~new_G556;
  assign new_G562 = ~new_G560 | ~new_G561;
  assign new_G586 = ~new_G553 | ~new_G554;
  assign new_G630 = new_G540 & new_G905;
  assign new_G634 = ~new_G540 | ~new_G905;
  assign new_G639 = ~new_G636;
  assign new_G642 = ~new_G3082 | ~new_G3085;
  assign new_G3086 = ~new_G3082;
  assign new_G644 = new_G460 & new_G636;
  assign new_G646 = ~new_G3098 | ~new_G3101;
  assign new_G3102 = ~new_G3098;
  assign new_G654 = ~G87 | ~new_G626;
  assign new_G660 = ~new_G657;
  assign new_G678 = ~new_G675;
  assign new_G804 = ~new_G860 | ~new_G776;
  assign new_G806 = ~new_G860 | ~new_G780;
  assign new_G855 = ~new_G736 | ~new_G707 | ~new_G721;
  assign new_G867 = ~new_G794 | ~new_G736 | ~new_G707 | ~new_G724;
  assign new_G903 = ~new_G3090 | ~new_G3093;
  assign new_G3094 = ~new_G3090;
  assign new_G912 = ~new_G3106 | ~new_G3109;
  assign new_G3110 = ~new_G3106;
  assign new_G915 = ~new_G861;
  assign new_G927 = ~new_G893;
  assign new_G941 = ~new_G864;
  assign new_G977 = new_G828 & new_G974;
  assign new_G978 = G150 & new_G975;
  assign new_G984 = new_G833 & new_G981;
  assign new_G985 = G159 & new_G982;
  assign new_G991 = G77 & new_G988;
  assign new_G992 = G50 & new_G989;
  assign new_G998 = new_G839 & new_G995;
  assign new_G999 = new_G828 & new_G996;
  assign new_G1005 = new_G845 & new_G1002;
  assign new_G1006 = new_G833 & new_G1003;
  assign new_G1012 = G107 & new_G1009;
  assign new_G1013 = G77 & new_G1010;
  assign new_G1019 = G116 & new_G1016;
  assign new_G1020 = new_G839 & new_G1017;
  assign new_G1026 = G283 & new_G1023;
  assign new_G1027 = new_G845 & new_G1024;
  assign new_G1060 = G200 & new_G1054;
  assign new_G1063 = new_G1048 & new_G1054;
  assign new_G1066 = new_G1049 & new_G1057;
  assign new_G1069 = new_G1050 & new_G1057;
  assign new_G1527 = ~new_G784 | ~new_G794;
  assign new_G1530 = ~new_G776 | ~new_G794;
  assign new_G1542 = ~new_G1541 | ~new_G707 | ~new_G721;
  assign new_G1563 = ~new_G784 | ~new_G724 | ~new_G732;
  assign new_G1572 = ~new_G724 | ~new_G784;
  assign new_G1581 = ~new_G1512;
  assign new_G1585 = ~new_G1512;
  assign new_G1589 = ~new_G1512;
  assign new_G1593 = ~new_G1512;
  assign new_G1597 = ~new_G1512;
  assign new_G1601 = ~new_G1512;
  assign new_G1605 = ~new_G1512;
  assign new_G1716 = ~new_G1681;
  assign new_G1718 = new_G1681 & new_G1699;
  assign new_G1723 = ~new_G1681;
  assign new_G1725 = new_G1681 & new_G1699;
  assign new_G1730 = ~new_G1681;
  assign new_G1732 = new_G1681 & new_G1699;
  assign new_G1737 = ~new_G1681;
  assign new_G1739 = new_G1681 & new_G1699;
  assign new_G1744 = ~new_G1681;
  assign new_G1746 = new_G1681 & new_G1699;
  assign new_G1751 = ~new_G1681;
  assign new_G1753 = new_G1681 & new_G1699;
  assign new_G1758 = ~new_G1681;
  assign new_G1760 = new_G1681 & new_G1699;
  assign new_G1765 = ~new_G1681;
  assign new_G1767 = new_G1681 & new_G1699;
  assign new_G1852 = new_G1834 & new_G1773;
  assign new_G1856 = ~G50 & ~new_G1773;
  assign new_G1870 = ~new_G807;
  assign new_G1902 = new_G1834 & new_G1773;
  assign new_G1906 = ~G58 & ~new_G1773;
  assign new_G1920 = ~new_G807;
  assign new_G1953 = new_G1834 & new_G1773;
  assign new_G1957 = ~G68 & ~new_G1773;
  assign new_G1971 = ~new_G807;
  assign new_G2003 = new_G1834 & new_G1773;
  assign new_G2007 = ~G77 & ~new_G1773;
  assign new_G2021 = ~new_G807;
  assign new_G2058 = new_G1834 & new_G1773;
  assign new_G2062 = ~G87 & ~new_G1773;
  assign new_G2076 = ~new_G823;
  assign new_G2110 = new_G1834 & new_G1773;
  assign new_G2114 = ~G97 & ~new_G1773;
  assign new_G2128 = ~new_G816;
  assign new_G2163 = new_G1834 & new_G1773;
  assign new_G2167 = ~G107 & ~new_G1773;
  assign new_G2181 = ~new_G816;
  assign new_G2215 = new_G1834 & new_G1773;
  assign new_G2219 = ~G116 & ~new_G1773;
  assign new_G2233 = ~new_G816;
  assign new_G2285 = new_G2278 & G213;
  assign new_G2288 = ~new_G2278 | ~G213;
  assign new_G2289 = G343 & new_G2278 & G213;
  assign new_G2293 = ~G343 | ~new_G2278 | ~G213;
  assign new_G2298 = G343 & new_G2278 & G213;
  assign new_G2302 = ~G343 | ~new_G2278 | ~G213;
  assign new_G2877 = new_G2874;
  assign new_G2983 = ~new_G2955 | ~new_G2956;
  assign new_G2986 = ~new_G2965 | ~new_G2966;
  assign new_G3014 = ~new_G3010;
  assign new_G3015 = ~new_G3010 | ~new_G3013;
  assign new_G3023 = ~new_G3017;
  assign new_G3024 = ~new_G3020;
  assign new_G3033 = ~new_G3027;
  assign new_G3034 = ~new_G3030;
  assign new_G3043 = ~new_G3037;
  assign new_G3044 = ~new_G3040;
  assign G355 = ~new_G354;
  assign new_G643 = ~new_G3079 | ~new_G3086;
  assign new_G647 = ~new_G3095 | ~new_G3102;
  assign new_G680 = new_G650 & new_G675;
  assign new_G904 = ~new_G3087 | ~new_G3094;
  assign new_G913 = ~new_G3103 | ~new_G3110;
  assign new_G920 = new_G588 & new_G915;
  assign new_G979 = new_G978 | new_G976 | new_G977;
  assign new_G993 = new_G992 | new_G990 | new_G991;
  assign new_G1000 = new_G999 | new_G997 | new_G998;
  assign new_G1007 = new_G1006 | new_G1004 | new_G1005;
  assign new_G1021 = new_G1020 | new_G1018 | new_G1019;
  assign new_G1028 = new_G1027 | new_G1025 | new_G1026;
  assign new_G1719 = G77 & new_G1716;
  assign new_G1721 = G223 & new_G1718;
  assign new_G1726 = G87 & new_G1723;
  assign new_G1728 = G226 & new_G1725;
  assign new_G1733 = G97 & new_G1730;
  assign new_G1735 = G232 & new_G1732;
  assign new_G1740 = G107 & new_G1737;
  assign new_G1742 = G238 & new_G1739;
  assign new_G1747 = G116 & new_G1744;
  assign new_G1749 = G244 & new_G1746;
  assign new_G1754 = G283 & new_G1751;
  assign new_G1756 = G250 & new_G1753;
  assign new_G1761 = G294 & new_G1758;
  assign new_G1763 = G257 & new_G1760;
  assign new_G1768 = G303 & new_G1765;
  assign new_G1770 = G264 & new_G1767;
  assign new_G1794 = new_G1791;
  assign new_G1799 = ~new_G1791;
  assign new_G1812 = new_G1809;
  assign new_G1817 = ~new_G1809;
  assign new_G1859 = new_G1852 & G50 & new_G1829;
  assign new_G1909 = new_G1902 & G58 & new_G1829;
  assign new_G1960 = new_G1953 & G68 & new_G1829;
  assign new_G2010 = new_G2003 & G77 & new_G1829;
  assign new_G2065 = new_G2058 & G87 & new_G2052;
  assign new_G2117 = new_G2110 & G97 & new_G2052;
  assign new_G2170 = new_G2163 & G107 & new_G2052;
  assign new_G2222 = new_G2215 & G116 & new_G2052;
  assign new_G2678 = ~new_G956;
  assign new_G2697 = ~new_G956;
  assign new_G2716 = ~new_G956;
  assign new_G2733 = ~new_G956;
  assign new_G2751 = ~new_G956;
  assign new_G2768 = ~new_G956;
  assign new_G2785 = ~new_G956;
  assign new_G2802 = ~new_G956;
  assign new_G3016 = ~new_G3007 | ~new_G3014;
  assign new_G3025 = ~new_G3020 | ~new_G3023;
  assign new_G3026 = ~new_G3017 | ~new_G3024;
  assign new_G3035 = ~new_G3030 | ~new_G3033;
  assign new_G3036 = ~new_G3027 | ~new_G3034;
  assign new_G3045 = ~new_G3040 | ~new_G3043;
  assign new_G3046 = ~new_G3037 | ~new_G3044;
  assign new_G2989 = ~new_G2983;
  assign new_G2990 = ~new_G2986;
  assign new_G610 = ~new_G804;
  assign new_G613 = new_G804 & new_G806;
  assign new_G616 = ~new_G806;
  assign new_G640 = ~new_G642 | ~new_G643;
  assign new_G648 = ~new_G646 | ~new_G647;
  assign new_G655 = G58 & new_G442 & new_G630 & new_G635;
  assign new_G665 = ~new_G804;
  assign new_G668 = new_G804 & new_G806;
  assign new_G671 = ~new_G806;
  assign new_G683 = ~new_G804;
  assign new_G685 = ~new_G806;
  assign new_G688 = new_G804 & new_G806;
  assign new_G694 = ~new_G804;
  assign new_G696 = ~new_G806;
  assign new_G699 = new_G804 & new_G806;
  assign new_G870 = new_G867;
  assign new_G887 = new_G867;
  assign new_G901 = ~new_G903 | ~new_G904;
  assign new_G910 = ~new_G912 | ~new_G913;
  assign new_G914 = ~new_G855;
  assign new_G916 = new_G855 & new_G861;
  assign new_G942 = ~new_G855;
  assign new_G943 = new_G864 & new_G855;
  assign new_G1072 = ~new_G1043 | ~new_G1069;
  assign new_G1084 = ~new_G1043 | ~new_G1066;
  assign new_G1096 = ~new_G1038 | ~new_G1069;
  assign new_G1108 = ~new_G1038 | ~new_G1066;
  assign new_G1120 = ~new_G1043 | ~new_G1063;
  assign new_G1132 = ~new_G1043 | ~new_G1060;
  assign new_G1144 = ~new_G1038 | ~new_G1063;
  assign new_G1156 = ~new_G1038 | ~new_G1060;
  assign new_G1533 = ~new_G1527;
  assign new_G1534 = ~new_G1530;
  assign new_G1535 = new_G1527 & new_G1530;
  assign new_G1545 = new_G1542;
  assign new_G1554 = new_G1542;
  assign new_G1610 = ~new_G1572;
  assign new_G1619 = ~new_G1572;
  assign new_G1628 = ~new_G1572;
  assign new_G1637 = ~new_G1572;
  assign new_G1646 = ~new_G1563;
  assign new_G1655 = ~new_G1563;
  assign new_G1664 = ~new_G1563;
  assign new_G1673 = ~new_G1563;
  assign new_G1722 = new_G1721 | new_G1719 | new_G1720;
  assign new_G1729 = new_G1728 | new_G1726 | new_G1727;
  assign new_G1736 = new_G1735 | new_G1733 | new_G1734;
  assign new_G1743 = new_G1742 | new_G1740 | new_G1741;
  assign new_G1750 = new_G1749 | new_G1747 | new_G1748;
  assign new_G1757 = new_G1756 | new_G1754 | new_G1755;
  assign new_G1764 = new_G1763 | new_G1761 | new_G1762;
  assign new_G1771 = new_G1770 | new_G1768 | new_G1769;
  assign new_G1853 = new_G979 & new_G1851;
  assign new_G1954 = new_G993 & new_G1952;
  assign new_G2004 = new_G1000 & new_G2002;
  assign new_G2059 = new_G1007 & new_G2057;
  assign new_G2164 = new_G1021 & new_G2162;
  assign new_G2216 = new_G1028 & new_G2214;
  assign new_G2485 = new_G2293;
  assign new_G2900 = new_G2877 & G2897;
  assign new_G2903 = ~new_G2877 | ~G2897;
  assign new_G2967 = new_G557;
  assign new_G2970 = new_G562;
  assign new_G2975 = new_G557;
  assign new_G2978 = new_G562;
  assign new_G3047 = ~new_G3015 | ~new_G3016;
  assign new_G3050 = ~new_G3025 | ~new_G3026;
  assign new_G3055 = ~new_G3035 | ~new_G3036;
  assign new_G3058 = ~new_G3045 | ~new_G3046;
  assign new_G574 = ~new_G2986 | ~new_G2989;
  assign new_G575 = ~new_G2983 | ~new_G2990;
  assign new_G617 = new_G501 & new_G613;
  assign new_G641 = new_G639 & new_G640 & new_G476;
  assign new_G649 = new_G530 & new_G648;
  assign new_G662 = new_G655 & new_G657;
  assign new_G672 = new_G513 & new_G668;
  assign new_G690 = new_G654 & new_G685;
  assign new_G691 = new_G540 & new_G688;
  assign new_G701 = new_G634 & new_G696;
  assign new_G702 = new_G526 & new_G699;
  assign new_G902 = ~new_G901;
  assign new_G911 = ~new_G910;
  assign new_G917 = new_G650 & new_G914;
  assign new_G923 = new_G586 & new_G916;
  assign new_G1538 = new_G442 & new_G1535;
  assign new_G1871 = new_G1870 & new_G1817 & G226;
  assign new_G1872 = new_G807 & new_G1817 & G274;
  assign new_G1873 = new_G1812 & new_G1722;
  assign new_G1921 = new_G1920 & new_G1817 & G232;
  assign new_G1922 = new_G807 & new_G1817 & G274;
  assign new_G1923 = new_G1812 & new_G1729;
  assign new_G1972 = new_G1971 & new_G1817 & G238;
  assign new_G1973 = new_G807 & new_G1817 & G274;
  assign new_G1974 = new_G1812 & new_G1736;
  assign new_G2022 = new_G2021 & new_G1817 & G244;
  assign new_G2023 = new_G807 & new_G1817 & G274;
  assign new_G2024 = new_G1812 & new_G1743;
  assign new_G2077 = new_G2076 & new_G1799 & G250;
  assign new_G2078 = new_G823 & new_G1799 & G274;
  assign new_G2079 = new_G1794 & new_G1750;
  assign new_G2129 = new_G2128 & new_G1799 & G257;
  assign new_G2130 = new_G816 & new_G1799 & G274;
  assign new_G2131 = new_G1794 & new_G1757;
  assign new_G2182 = new_G2181 & new_G1799 & G264;
  assign new_G2183 = new_G816 & new_G1799 & G274;
  assign new_G2184 = new_G1794 & new_G1764;
  assign new_G2234 = new_G2233 & new_G1799 & G270;
  assign new_G2235 = new_G816 & new_G1799 & G274;
  assign new_G2236 = new_G1794 & new_G1771;
  assign new_G2973 = ~new_G2967;
  assign new_G2974 = ~new_G2970;
  assign new_G2981 = ~new_G2975;
  assign new_G2982 = ~new_G2978;
  assign new_G576 = ~new_G574 | ~new_G575;
  assign new_G3053 = ~new_G3047;
  assign new_G3054 = ~new_G3050;
  assign new_G3061 = ~new_G3055;
  assign new_G3062 = ~new_G3058;
  assign new_G645 = new_G641 | new_G644;
  assign new_G926 = ~new_G887;
  assign new_G928 = new_G887 & new_G893;
  assign new_G947 = new_G649 & new_G942;
  assign new_G983 = new_G902 & new_G980;
  assign new_G1011 = new_G911 & new_G1008;
  assign new_G1075 = new_G1072;
  assign new_G1087 = new_G1084;
  assign new_G1099 = new_G1096;
  assign new_G1111 = new_G1108;
  assign new_G1123 = new_G1120;
  assign new_G1135 = new_G1132;
  assign new_G1147 = new_G1144;
  assign new_G1159 = new_G1156;
  assign new_G1168 = new_G1072;
  assign new_G1177 = new_G1084;
  assign new_G1186 = new_G1096;
  assign new_G1195 = new_G1108;
  assign new_G1204 = new_G1120;
  assign new_G1213 = new_G1132;
  assign new_G1222 = new_G1144;
  assign new_G1231 = new_G1156;
  assign new_G1609 = ~new_G1545;
  assign new_G1611 = new_G1545 & new_G1572;
  assign new_G1618 = ~new_G1545;
  assign new_G1620 = new_G1545 & new_G1572;
  assign new_G1627 = ~new_G1545;
  assign new_G1629 = new_G1545 & new_G1572;
  assign new_G1636 = ~new_G1545;
  assign new_G1638 = new_G1545 & new_G1572;
  assign new_G1645 = ~new_G1554;
  assign new_G1647 = new_G1554 & new_G1563;
  assign new_G1654 = ~new_G1554;
  assign new_G1656 = new_G1554 & new_G1563;
  assign new_G1663 = ~new_G1554;
  assign new_G1665 = new_G1554 & new_G1563;
  assign new_G1672 = ~new_G1554;
  assign new_G1674 = new_G1554 & new_G1563;
  assign new_G1862 = new_G1859 | new_G1853 | new_G1856;
  assign new_G1866 = ~new_G1859 & ~new_G1853 & ~new_G1856;
  assign new_G1874 = new_G1873 | new_G1871 | new_G1872;
  assign new_G1924 = new_G1923 | new_G1921 | new_G1922;
  assign new_G1963 = new_G1960 | new_G1954 | new_G1957;
  assign new_G1967 = ~new_G1960 & ~new_G1954 & ~new_G1957;
  assign new_G1975 = new_G1974 | new_G1972 | new_G1973;
  assign new_G2013 = new_G2010 | new_G2004 | new_G2007;
  assign new_G2017 = ~new_G2010 & ~new_G2004 & ~new_G2007;
  assign new_G2025 = new_G2024 | new_G2022 | new_G2023;
  assign new_G2068 = new_G2065 | new_G2059 | new_G2062;
  assign new_G2072 = ~new_G2065 & ~new_G2059 & ~new_G2062;
  assign new_G2080 = new_G2079 | new_G2077 | new_G2078;
  assign new_G2132 = new_G2131 | new_G2129 | new_G2130;
  assign new_G2173 = new_G2170 | new_G2164 | new_G2167;
  assign new_G2177 = ~new_G2170 & ~new_G2164 & ~new_G2167;
  assign new_G2185 = new_G2184 | new_G2182 | new_G2183;
  assign new_G2225 = new_G2222 | new_G2216 | new_G2219;
  assign new_G2229 = ~new_G2222 & ~new_G2216 & ~new_G2219;
  assign new_G2237 = new_G2236 | new_G2234 | new_G2235;
  assign new_G2488 = ~new_G2485;
  assign new_G2679 = ~new_G870;
  assign new_G2680 = new_G956 & new_G870;
  assign new_G2698 = ~new_G870;
  assign new_G2699 = new_G956 & new_G870;
  assign new_G2717 = ~new_G870;
  assign new_G2718 = new_G956 & new_G870;
  assign new_G2734 = ~new_G870;
  assign new_G2735 = new_G956 & new_G870;
  assign new_G2752 = ~new_G870;
  assign new_G2753 = new_G956 & new_G870;
  assign new_G2769 = ~new_G870;
  assign new_G2770 = new_G956 & new_G870;
  assign new_G2786 = ~new_G870;
  assign new_G2787 = new_G956 & new_G870;
  assign new_G2803 = ~new_G870;
  assign new_G2804 = new_G956 & new_G870;
  assign new_G359 = new_G923 | new_G917 | new_G920;
  assign new_G1029 = ~new_G923 & ~new_G917 & ~new_G920;
  assign new_G565 = ~new_G2970 | ~new_G2973;
  assign new_G566 = ~new_G2967 | ~new_G2974;
  assign new_G569 = ~new_G2978 | ~new_G2981;
  assign new_G570 = ~new_G2975 | ~new_G2982;
  assign new_G589 = ~new_G3050 | ~new_G3053;
  assign new_G590 = ~new_G3047 | ~new_G3054;
  assign new_G595 = ~new_G3058 | ~new_G3061;
  assign new_G596 = ~new_G3055 | ~new_G3062;
  assign new_G929 = new_G650 & new_G926;
  assign new_G938 = new_G630 & new_G928;
  assign new_G944 = new_G645 & new_G941;
  assign new_G986 = new_G985 | new_G983 | new_G984;
  assign new_G1014 = new_G1013 | new_G1011 | new_G1012;
  assign new_G1616 = new_G442 & new_G1611;
  assign new_G1625 = new_G456 & new_G1620;
  assign new_G1634 = new_G463 & new_G1629;
  assign new_G1643 = new_G479 & new_G1638;
  assign new_G360 = ~new_G1029;
  assign new_G567 = ~new_G565 | ~new_G566;
  assign new_G571 = ~new_G569 | ~new_G570;
  assign new_G579 = new_G576;
  assign new_G591 = ~new_G589 | ~new_G590;
  assign new_G597 = ~new_G595 | ~new_G596;
  assign new_G614 = new_G576 & new_G610;
  assign new_G1240 = ~new_G1075;
  assign new_G1241 = ~new_G1087;
  assign new_G1242 = ~new_G1099;
  assign new_G1243 = ~new_G1111;
  assign new_G1244 = ~new_G1123;
  assign new_G1245 = ~new_G1135;
  assign new_G1246 = ~new_G1147;
  assign new_G1247 = ~new_G1159;
  assign new_G1257 = ~new_G1075;
  assign new_G1258 = ~new_G1087;
  assign new_G1259 = ~new_G1099;
  assign new_G1260 = ~new_G1111;
  assign new_G1261 = ~new_G1123;
  assign new_G1262 = ~new_G1135;
  assign new_G1263 = ~new_G1147;
  assign new_G1264 = ~new_G1159;
  assign new_G1274 = ~new_G1075;
  assign new_G1275 = ~new_G1087;
  assign new_G1276 = ~new_G1099;
  assign new_G1277 = ~new_G1111;
  assign new_G1278 = ~new_G1123;
  assign new_G1279 = ~new_G1135;
  assign new_G1280 = ~new_G1147;
  assign new_G1281 = ~new_G1159;
  assign new_G1291 = ~new_G1075;
  assign new_G1292 = ~new_G1087;
  assign new_G1293 = ~new_G1099;
  assign new_G1294 = ~new_G1111;
  assign new_G1295 = ~new_G1123;
  assign new_G1296 = ~new_G1135;
  assign new_G1297 = ~new_G1147;
  assign new_G1298 = ~new_G1159;
  assign new_G1308 = ~new_G1075;
  assign new_G1309 = ~new_G1087;
  assign new_G1310 = ~new_G1099;
  assign new_G1311 = ~new_G1111;
  assign new_G1312 = ~new_G1123;
  assign new_G1313 = ~new_G1135;
  assign new_G1314 = ~new_G1147;
  assign new_G1315 = ~new_G1159;
  assign new_G1325 = ~new_G1075;
  assign new_G1326 = ~new_G1087;
  assign new_G1327 = ~new_G1099;
  assign new_G1328 = ~new_G1111;
  assign new_G1329 = ~new_G1123;
  assign new_G1330 = ~new_G1135;
  assign new_G1331 = ~new_G1147;
  assign new_G1332 = ~new_G1159;
  assign new_G1342 = ~new_G1075;
  assign new_G1343 = ~new_G1087;
  assign new_G1344 = ~new_G1099;
  assign new_G1345 = ~new_G1111;
  assign new_G1346 = ~new_G1123;
  assign new_G1347 = ~new_G1135;
  assign new_G1348 = ~new_G1147;
  assign new_G1349 = ~new_G1159;
  assign new_G1359 = ~new_G1075;
  assign new_G1360 = ~new_G1087;
  assign new_G1361 = ~new_G1099;
  assign new_G1362 = ~new_G1111;
  assign new_G1363 = ~new_G1123;
  assign new_G1364 = ~new_G1135;
  assign new_G1365 = ~new_G1147;
  assign new_G1366 = ~new_G1159;
  assign new_G1376 = ~new_G1168;
  assign new_G1377 = ~new_G1177;
  assign new_G1378 = ~new_G1186;
  assign new_G1379 = ~new_G1195;
  assign new_G1380 = ~new_G1204;
  assign new_G1381 = ~new_G1213;
  assign new_G1382 = ~new_G1222;
  assign new_G1383 = ~new_G1231;
  assign new_G1393 = ~new_G1168;
  assign new_G1394 = ~new_G1177;
  assign new_G1395 = ~new_G1186;
  assign new_G1396 = ~new_G1195;
  assign new_G1397 = ~new_G1204;
  assign new_G1398 = ~new_G1213;
  assign new_G1399 = ~new_G1222;
  assign new_G1400 = ~new_G1231;
  assign new_G1410 = ~new_G1168;
  assign new_G1411 = ~new_G1177;
  assign new_G1412 = ~new_G1186;
  assign new_G1413 = ~new_G1195;
  assign new_G1414 = ~new_G1204;
  assign new_G1415 = ~new_G1213;
  assign new_G1416 = ~new_G1222;
  assign new_G1417 = ~new_G1231;
  assign new_G1427 = ~new_G1168;
  assign new_G1428 = ~new_G1177;
  assign new_G1429 = ~new_G1186;
  assign new_G1430 = ~new_G1195;
  assign new_G1431 = ~new_G1204;
  assign new_G1432 = ~new_G1213;
  assign new_G1433 = ~new_G1222;
  assign new_G1434 = ~new_G1231;
  assign new_G1444 = ~new_G1168;
  assign new_G1445 = ~new_G1177;
  assign new_G1446 = ~new_G1186;
  assign new_G1447 = ~new_G1195;
  assign new_G1448 = ~new_G1204;
  assign new_G1449 = ~new_G1213;
  assign new_G1450 = ~new_G1222;
  assign new_G1451 = ~new_G1231;
  assign new_G1461 = ~new_G1168;
  assign new_G1462 = ~new_G1177;
  assign new_G1463 = ~new_G1186;
  assign new_G1464 = ~new_G1195;
  assign new_G1465 = ~new_G1204;
  assign new_G1466 = ~new_G1213;
  assign new_G1467 = ~new_G1222;
  assign new_G1468 = ~new_G1231;
  assign new_G1478 = ~new_G1168;
  assign new_G1479 = ~new_G1177;
  assign new_G1480 = ~new_G1186;
  assign new_G1481 = ~new_G1195;
  assign new_G1482 = ~new_G1204;
  assign new_G1483 = ~new_G1213;
  assign new_G1484 = ~new_G1222;
  assign new_G1485 = ~new_G1231;
  assign new_G1495 = ~new_G1168;
  assign new_G1496 = ~new_G1177;
  assign new_G1497 = ~new_G1186;
  assign new_G1498 = ~new_G1195;
  assign new_G1499 = ~new_G1204;
  assign new_G1500 = ~new_G1213;
  assign new_G1501 = ~new_G1222;
  assign new_G1502 = ~new_G1231;
  assign new_G1877 = new_G1874;
  assign new_G1880 = ~new_G1874;
  assign new_G1891 = ~new_G1866;
  assign new_G1903 = new_G986 & new_G1901;
  assign new_G1927 = new_G1924;
  assign new_G1930 = ~new_G1924;
  assign new_G1978 = new_G1975;
  assign new_G1981 = ~new_G1975;
  assign new_G1992 = ~new_G1967;
  assign new_G2028 = new_G2025;
  assign new_G2031 = ~new_G2025;
  assign new_G2042 = ~new_G2017;
  assign new_G2085 = new_G2080;
  assign new_G2088 = ~new_G2080;
  assign new_G2099 = ~new_G2072;
  assign new_G2111 = new_G1014 & new_G2109;
  assign new_G2137 = new_G2132;
  assign new_G2140 = ~new_G2132;
  assign new_G2190 = new_G2185;
  assign new_G2193 = ~new_G2185;
  assign new_G2204 = ~new_G2177;
  assign new_G2242 = new_G2237;
  assign new_G2245 = ~new_G2237;
  assign new_G2256 = ~new_G2229;
  assign new_G2320 = new_G2285 & new_G1862;
  assign new_G2341 = new_G2289 & new_G1963;
  assign new_G2354 = new_G2289 & new_G2013;
  assign new_G2367 = new_G2289 & new_G2068;
  assign new_G2383 = new_G2298 & new_G2173;
  assign new_G2391 = new_G2298 & new_G2225;
  assign new_G2474 = ~new_G2080;
  assign new_G2475 = ~new_G2132;
  assign new_G2476 = ~new_G2185;
  assign new_G2477 = ~new_G2237;
  assign new_G2482 = new_G2481 & new_G2237 & new_G2185 & new_G2080 & new_G2132;
  assign G361 = ~new_G359 | ~new_G360;
  assign new_G568 = ~new_G567;
  assign new_G618 = new_G617 | new_G614 | new_G616;
  assign new_G1248 = G124 & new_G1240;
  assign new_G1249 = G159 & new_G1241;
  assign new_G1250 = G150 & new_G1242;
  assign new_G1251 = G143 & new_G1243;
  assign new_G1252 = G137 & new_G1244;
  assign new_G1253 = G132 & new_G1245;
  assign new_G1254 = G128 & new_G1246;
  assign new_G1255 = G125 & new_G1247;
  assign new_G1265 = G125 & new_G1257;
  assign new_G1266 = new_G432 & new_G1258;
  assign new_G1267 = G159 & new_G1259;
  assign new_G1268 = G150 & new_G1260;
  assign new_G1269 = G143 & new_G1261;
  assign new_G1270 = G137 & new_G1262;
  assign new_G1271 = G132 & new_G1263;
  assign new_G1272 = G128 & new_G1264;
  assign new_G1282 = G128 & new_G1274;
  assign new_G1283 = new_G447 & new_G1275;
  assign new_G1284 = new_G432 & new_G1276;
  assign new_G1285 = G159 & new_G1277;
  assign new_G1286 = G150 & new_G1278;
  assign new_G1287 = G143 & new_G1279;
  assign new_G1288 = G137 & new_G1280;
  assign new_G1289 = G132 & new_G1281;
  assign new_G1299 = G132 & new_G1291;
  assign new_G1300 = new_G467 & new_G1292;
  assign new_G1301 = new_G447 & new_G1293;
  assign new_G1302 = new_G432 & new_G1294;
  assign new_G1303 = G159 & new_G1295;
  assign new_G1304 = G150 & new_G1296;
  assign new_G1305 = G143 & new_G1297;
  assign new_G1306 = G137 & new_G1298;
  assign new_G1316 = G137 & new_G1308;
  assign new_G1317 = new_G483 & new_G1309;
  assign new_G1318 = new_G467 & new_G1310;
  assign new_G1319 = new_G447 & new_G1311;
  assign new_G1320 = new_G432 & new_G1312;
  assign new_G1321 = G159 & new_G1313;
  assign new_G1322 = G150 & new_G1314;
  assign new_G1323 = G143 & new_G1315;
  assign new_G1333 = G143 & new_G1325;
  assign new_G1334 = new_G492 & new_G1326;
  assign new_G1335 = new_G483 & new_G1327;
  assign new_G1336 = new_G467 & new_G1328;
  assign new_G1337 = new_G447 & new_G1329;
  assign new_G1338 = new_G432 & new_G1330;
  assign new_G1339 = G159 & new_G1331;
  assign new_G1340 = G150 & new_G1332;
  assign new_G1350 = G150 & new_G1342;
  assign new_G1351 = new_G504 & new_G1343;
  assign new_G1352 = new_G492 & new_G1344;
  assign new_G1353 = new_G483 & new_G1345;
  assign new_G1354 = new_G467 & new_G1346;
  assign new_G1355 = new_G447 & new_G1347;
  assign new_G1356 = new_G432 & new_G1348;
  assign new_G1357 = G159 & new_G1349;
  assign new_G1367 = G159 & new_G1359;
  assign new_G1368 = new_G517 & new_G1360;
  assign new_G1369 = new_G504 & new_G1361;
  assign new_G1370 = new_G492 & new_G1362;
  assign new_G1371 = new_G483 & new_G1363;
  assign new_G1372 = new_G467 & new_G1364;
  assign new_G1373 = new_G447 & new_G1365;
  assign new_G1374 = new_G432 & new_G1366;
  assign new_G1384 = G283 & new_G1376;
  assign new_G1385 = new_G447 & new_G1377;
  assign new_G1386 = new_G467 & new_G1378;
  assign new_G1387 = new_G483 & new_G1379;
  assign new_G1388 = new_G492 & new_G1380;
  assign new_G1389 = new_G504 & new_G1381;
  assign new_G1390 = new_G517 & new_G1382;
  assign new_G1391 = new_G530 & new_G1383;
  assign new_G1401 = G294 & new_G1393;
  assign new_G1402 = new_G467 & new_G1394;
  assign new_G1403 = new_G483 & new_G1395;
  assign new_G1404 = new_G492 & new_G1396;
  assign new_G1405 = new_G504 & new_G1397;
  assign new_G1406 = new_G517 & new_G1398;
  assign new_G1407 = new_G530 & new_G1399;
  assign new_G1408 = G283 & new_G1400;
  assign new_G1418 = G303 & new_G1410;
  assign new_G1419 = new_G483 & new_G1411;
  assign new_G1420 = new_G492 & new_G1412;
  assign new_G1421 = new_G504 & new_G1413;
  assign new_G1422 = new_G517 & new_G1414;
  assign new_G1423 = new_G530 & new_G1415;
  assign new_G1424 = G283 & new_G1416;
  assign new_G1425 = G294 & new_G1417;
  assign new_G1435 = G311 & new_G1427;
  assign new_G1436 = new_G492 & new_G1428;
  assign new_G1437 = new_G504 & new_G1429;
  assign new_G1438 = new_G517 & new_G1430;
  assign new_G1439 = new_G530 & new_G1431;
  assign new_G1440 = G283 & new_G1432;
  assign new_G1441 = G294 & new_G1433;
  assign new_G1442 = G303 & new_G1434;
  assign new_G1452 = G317 & new_G1444;
  assign new_G1453 = new_G504 & new_G1445;
  assign new_G1454 = new_G517 & new_G1446;
  assign new_G1455 = new_G530 & new_G1447;
  assign new_G1456 = G283 & new_G1448;
  assign new_G1457 = G294 & new_G1449;
  assign new_G1458 = G303 & new_G1450;
  assign new_G1459 = G311 & new_G1451;
  assign new_G1469 = G322 & new_G1461;
  assign new_G1470 = new_G517 & new_G1462;
  assign new_G1471 = new_G530 & new_G1463;
  assign new_G1472 = G283 & new_G1464;
  assign new_G1473 = G294 & new_G1465;
  assign new_G1474 = G303 & new_G1466;
  assign new_G1475 = G311 & new_G1467;
  assign new_G1476 = G317 & new_G1468;
  assign new_G1486 = G326 & new_G1478;
  assign new_G1487 = new_G530 & new_G1479;
  assign new_G1488 = G283 & new_G1480;
  assign new_G1489 = G294 & new_G1481;
  assign new_G1490 = G303 & new_G1482;
  assign new_G1491 = G311 & new_G1483;
  assign new_G1492 = G317 & new_G1484;
  assign new_G1493 = G322 & new_G1485;
  assign new_G1503 = G329 & new_G1495;
  assign new_G1504 = G283 & new_G1496;
  assign new_G1505 = G294 & new_G1497;
  assign new_G1506 = G303 & new_G1498;
  assign new_G1507 = G311 & new_G1499;
  assign new_G1508 = G317 & new_G1500;
  assign new_G1509 = G322 & new_G1501;
  assign new_G1510 = G326 & new_G1502;
  assign new_G2483 = new_G2478 & new_G2477 & new_G2476 & new_G2474 & new_G2475;
  assign new_G600 = new_G597;
  assign new_G661 = new_G568 & new_G660;
  assign new_G669 = new_G597 & new_G665;
  assign new_G679 = new_G591 & new_G678;
  assign new_G1256 = ~new_G1255 & ~new_G1254 & ~new_G1253 & ~new_G1252 & ~new_G1251 & ~new_G1250 & ~new_G1248 & ~new_G1249;
  assign new_G1273 = ~new_G1272 & ~new_G1271 & ~new_G1270 & ~new_G1269 & ~new_G1268 & ~new_G1267 & ~new_G1265 & ~new_G1266;
  assign new_G1290 = ~new_G1289 & ~new_G1288 & ~new_G1287 & ~new_G1286 & ~new_G1285 & ~new_G1284 & ~new_G1282 & ~new_G1283;
  assign new_G1307 = ~new_G1306 & ~new_G1305 & ~new_G1304 & ~new_G1303 & ~new_G1302 & ~new_G1301 & ~new_G1299 & ~new_G1300;
  assign new_G1324 = ~new_G1323 & ~new_G1322 & ~new_G1321 & ~new_G1320 & ~new_G1319 & ~new_G1318 & ~new_G1316 & ~new_G1317;
  assign new_G1341 = ~new_G1340 & ~new_G1339 & ~new_G1338 & ~new_G1337 & ~new_G1336 & ~new_G1335 & ~new_G1333 & ~new_G1334;
  assign new_G1358 = ~new_G1357 & ~new_G1356 & ~new_G1355 & ~new_G1354 & ~new_G1353 & ~new_G1352 & ~new_G1350 & ~new_G1351;
  assign new_G1375 = ~new_G1374 & ~new_G1373 & ~new_G1372 & ~new_G1371 & ~new_G1370 & ~new_G1369 & ~new_G1367 & ~new_G1368;
  assign new_G1392 = ~new_G1391 & ~new_G1390 & ~new_G1389 & ~new_G1388 & ~new_G1387 & ~new_G1386 & ~new_G1384 & ~new_G1385;
  assign new_G1409 = ~new_G1408 & ~new_G1407 & ~new_G1406 & ~new_G1405 & ~new_G1404 & ~new_G1403 & ~new_G1401 & ~new_G1402;
  assign new_G1426 = ~new_G1425 & ~new_G1424 & ~new_G1423 & ~new_G1422 & ~new_G1421 & ~new_G1420 & ~new_G1418 & ~new_G1419;
  assign new_G1443 = ~new_G1442 & ~new_G1441 & ~new_G1440 & ~new_G1439 & ~new_G1438 & ~new_G1437 & ~new_G1435 & ~new_G1436;
  assign new_G1460 = ~new_G1459 & ~new_G1458 & ~new_G1457 & ~new_G1456 & ~new_G1455 & ~new_G1454 & ~new_G1452 & ~new_G1453;
  assign new_G1477 = ~new_G1476 & ~new_G1475 & ~new_G1474 & ~new_G1473 & ~new_G1472 & ~new_G1471 & ~new_G1469 & ~new_G1470;
  assign new_G1494 = ~new_G1493 & ~new_G1492 & ~new_G1491 & ~new_G1490 & ~new_G1489 & ~new_G1488 & ~new_G1486 & ~new_G1487;
  assign new_G1511 = ~new_G1510 & ~new_G1509 & ~new_G1508 & ~new_G1507 & ~new_G1506 & ~new_G1505 & ~new_G1503 & ~new_G1504;
  assign new_G1652 = new_G618 & new_G1647;
  assign new_G1883 = new_G1877 & G169 & new_G1862;
  assign new_G1886 = new_G1880 & G179 & new_G1862;
  assign new_G1889 = new_G1880 & G190 & new_G1866;
  assign new_G1890 = new_G1877 & G200 & new_G1866;
  assign new_G1912 = new_G1909 | new_G1903 | new_G1906;
  assign new_G1916 = ~new_G1909 & ~new_G1903 & ~new_G1906;
  assign new_G1984 = new_G1978 & G169 & new_G1963;
  assign new_G1987 = new_G1981 & G179 & new_G1963;
  assign new_G1990 = new_G1981 & G190 & new_G1967;
  assign new_G1991 = new_G1978 & G200 & new_G1967;
  assign new_G2034 = new_G2028 & G169 & new_G2013;
  assign new_G2037 = new_G2031 & G179 & new_G2013;
  assign new_G2040 = new_G2031 & G190 & new_G2017;
  assign new_G2041 = new_G2028 & G200 & new_G2017;
  assign new_G2091 = new_G2085 & G169 & new_G2068;
  assign new_G2094 = new_G2088 & G179 & new_G2068;
  assign new_G2097 = new_G2088 & G190 & new_G2072;
  assign new_G2098 = new_G2085 & G200 & new_G2072;
  assign new_G2120 = new_G2117 | new_G2111 | new_G2114;
  assign new_G2124 = ~new_G2117 & ~new_G2111 & ~new_G2114;
  assign new_G2196 = new_G2190 & G169 & new_G2173;
  assign new_G2199 = new_G2193 & G179 & new_G2173;
  assign new_G2202 = new_G2193 & G190 & new_G2177;
  assign new_G2203 = new_G2190 & G200 & new_G2177;
  assign new_G2248 = new_G2242 & G169 & new_G2225;
  assign new_G2251 = new_G2245 & G179 & new_G2225;
  assign new_G2254 = new_G2245 & G190 & new_G2229;
  assign new_G2255 = new_G2242 & G200 & new_G2229;
  assign new_G2484 = new_G2482 | new_G2483;
  assign new_G2991 = new_G571;
  assign new_G2994 = new_G579;
  assign new_G2999 = new_G571;
  assign new_G3002 = new_G579;
  assign new_G3063 = new_G591;
  assign new_G3071 = new_G591;
  assign new_G3124 = new_G2320;
  assign new_G3134 = new_G2320;
  assign new_G3158 = new_G2341;
  assign new_G3166 = new_G2341;
  assign new_G3174 = new_G2354;
  assign new_G3182 = new_G2354;
  assign new_G3190 = new_G2367;
  assign new_G3200 = new_G2367;
  assign new_G3224 = new_G2383;
  assign new_G3232 = new_G2383;
  assign new_G3240 = new_G2391;
  assign new_G3248 = new_G2391;
  assign new_G663 = ~new_G661 & ~new_G662;
  assign new_G673 = new_G672 | new_G669 | new_G671;
  assign new_G681 = ~new_G679 & ~new_G680;
  assign new_G1536 = new_G1256 & new_G1533;
  assign new_G1537 = new_G1392 & new_G1534;
  assign new_G1582 = new_G1273 & new_G1581;
  assign new_G1583 = new_G1409 & new_G1512;
  assign new_G1586 = new_G1290 & new_G1585;
  assign new_G1587 = new_G1426 & new_G1512;
  assign new_G1590 = new_G1307 & new_G1589;
  assign new_G1591 = new_G1443 & new_G1512;
  assign new_G1594 = new_G1324 & new_G1593;
  assign new_G1595 = new_G1460 & new_G1512;
  assign new_G1598 = new_G1341 & new_G1597;
  assign new_G1599 = new_G1477 & new_G1512;
  assign new_G1602 = new_G1358 & new_G1601;
  assign new_G1603 = new_G1494 & new_G1512;
  assign new_G1606 = new_G1375 & new_G1605;
  assign new_G1607 = new_G1511 & new_G1512;
  assign new_G1894 = new_G1891 | new_G1889 | new_G1890;
  assign new_G1997 = new_G1992 | new_G1990 | new_G1991;
  assign new_G2047 = new_G2042 | new_G2040 | new_G2041;
  assign new_G2102 = new_G2099 | new_G2097 | new_G2098;
  assign new_G2209 = new_G2204 | new_G2202 | new_G2203;
  assign new_G2261 = new_G2256 | new_G2254 | new_G2255;
  assign new_G2489 = new_G2484 & new_G2488;
  assign new_G3005 = ~new_G2999;
  assign new_G3006 = ~new_G3002;
  assign new_G3077 = ~new_G3071;
  assign new_G3069 = ~new_G3063;
  assign new_G2997 = ~new_G2991;
  assign new_G2998 = ~new_G2994;
  assign new_G689 = new_G681 & new_G683;
  assign new_G700 = new_G663 & new_G694;
  assign new_G1539 = new_G1538 | new_G1536 | new_G1537;
  assign new_G1584 = new_G1582 | new_G1583;
  assign new_G1588 = new_G1586 | new_G1587;
  assign new_G1592 = new_G1590 | new_G1591;
  assign new_G1596 = new_G1594 | new_G1595;
  assign new_G1600 = new_G1598 | new_G1599;
  assign new_G1604 = new_G1602 | new_G1603;
  assign new_G1608 = new_G1606 | new_G1607;
  assign new_G1661 = new_G673 & new_G1656;
  assign new_G1892 = new_G1883 | new_G1886;
  assign new_G1893 = ~new_G1883 & ~new_G1886;
  assign new_G1933 = new_G1927 & G169 & new_G1912;
  assign new_G1936 = new_G1930 & G179 & new_G1912;
  assign new_G1939 = new_G1930 & G190 & new_G1916;
  assign new_G1940 = new_G1927 & G200 & new_G1916;
  assign new_G1941 = ~new_G1916;
  assign new_G1993 = new_G1984 | new_G1987;
  assign new_G1996 = ~new_G1984 & ~new_G1987;
  assign new_G2043 = new_G2034 | new_G2037;
  assign new_G2046 = ~new_G2034 & ~new_G2037;
  assign new_G2100 = new_G2091 | new_G2094;
  assign new_G2101 = ~new_G2091 & ~new_G2094;
  assign new_G2143 = new_G2137 & G169 & new_G2120;
  assign new_G2146 = new_G2140 & G179 & new_G2120;
  assign new_G2149 = new_G2140 & G190 & new_G2124;
  assign new_G2150 = new_G2137 & G200 & new_G2124;
  assign new_G2151 = ~new_G2124;
  assign new_G2205 = new_G2196 | new_G2199;
  assign new_G2208 = ~new_G2196 & ~new_G2199;
  assign new_G2257 = new_G2248 | new_G2251;
  assign new_G2260 = ~new_G2248 & ~new_G2251;
  assign new_G3138 = ~new_G3134;
  assign new_G2328 = new_G2285 & new_G1912;
  assign new_G3162 = ~new_G3158;
  assign new_G3170 = ~new_G3166;
  assign new_G3178 = ~new_G3174;
  assign new_G3186 = ~new_G3182;
  assign new_G3204 = ~new_G3200;
  assign new_G2375 = new_G2298 & new_G2120;
  assign new_G3236 = ~new_G3232;
  assign new_G3244 = ~new_G3240;
  assign new_G3252 = ~new_G3248;
  assign new_G3228 = ~new_G3224;
  assign new_G3066 = new_G600;
  assign new_G3074 = new_G600;
  assign new_G3128 = ~new_G3124;
  assign new_G3194 = ~new_G3190;
  assign new_G619 = ~new_G2994 | ~new_G2997;
  assign new_G620 = ~new_G2991 | ~new_G2998;
  assign new_G582 = ~new_G3002 | ~new_G3005;
  assign new_G583 = ~new_G2999 | ~new_G3006;
  assign new_G692 = new_G691 | new_G689 | new_G690;
  assign new_G703 = new_G702 | new_G700 | new_G701;
  assign new_G1612 = new_G1539 & new_G1609;
  assign new_G1621 = new_G1584 & new_G1618;
  assign new_G1630 = new_G1588 & new_G1627;
  assign new_G1639 = new_G1592 & new_G1636;
  assign new_G1648 = new_G1596 & new_G1645;
  assign new_G1657 = new_G1600 & new_G1654;
  assign new_G1666 = new_G1604 & new_G1663;
  assign new_G1675 = new_G1608 & new_G1672;
  assign new_G1895 = new_G1893 & new_G1894;
  assign new_G1946 = new_G1941 | new_G1939 | new_G1940;
  assign new_G1998 = new_G1996 & new_G1997;
  assign new_G2048 = new_G2046 & new_G2047;
  assign new_G2103 = new_G2101 & new_G2102;
  assign new_G2156 = new_G2151 | new_G2149 | new_G2150;
  assign new_G2210 = new_G2208 & new_G2209;
  assign new_G2262 = new_G2260 & new_G2261;
  assign new_G2271 = ~new_G1892;
  assign new_G2311 = ~new_G2100;
  assign new_G356 = ~new_G619 | ~new_G620;
  assign new_G357 = ~new_G582 | ~new_G583;
  assign new_G603 = ~new_G3074 | ~new_G3077;
  assign new_G3078 = ~new_G3074;
  assign new_G606 = ~new_G3066 | ~new_G3069;
  assign new_G3070 = ~new_G3066;
  assign new_G1670 = new_G703 & new_G1665;
  assign new_G1679 = new_G692 & new_G1674;
  assign new_G1942 = new_G1933 | new_G1936;
  assign new_G1945 = ~new_G1933 & ~new_G1936;
  assign new_G2152 = new_G2143 | new_G2146;
  assign new_G2155 = ~new_G2143 & ~new_G2146;
  assign new_G2445 = new_G1993 & new_G2293;
  assign new_G2448 = new_G2043 & new_G2293;
  assign new_G2455 = new_G2205 & new_G2302;
  assign new_G2458 = new_G2257 & new_G2302;
  assign new_G3142 = new_G2328;
  assign new_G3150 = new_G2328;
  assign new_G3208 = new_G2375;
  assign new_G3216 = new_G2375;
  assign G358 = ~new_G356 | ~new_G357;
  assign new_G604 = ~new_G3071 | ~new_G3078;
  assign new_G607 = ~new_G3063 | ~new_G3070;
  assign new_G1947 = new_G1945 & new_G1946;
  assign new_G2157 = new_G2155 & new_G2156;
  assign new_G2317 = new_G1895;
  assign new_G2338 = new_G1998;
  assign new_G2351 = new_G2048;
  assign new_G2364 = new_G2103;
  assign new_G2380 = new_G2210;
  assign new_G2388 = new_G2262;
  assign new_G605 = ~new_G603 | ~new_G604;
  assign new_G608 = ~new_G606 | ~new_G607;
  assign new_G2272 = ~new_G1895 | ~new_G1942;
  assign new_G2312 = ~new_G2103 | ~new_G2152;
  assign new_G3146 = ~new_G3142;
  assign new_G3154 = ~new_G3150;
  assign new_G3220 = ~new_G3216;
  assign new_G3212 = ~new_G3208;
  assign new_G2444 = new_G1942 & new_G2288;
  assign new_G2451 = new_G2448;
  assign new_G2454 = new_G2152 & new_G2293;
  assign new_G2461 = new_G2458;
  assign new_G2530 = ~new_G2445;
  assign new_G3323 = new_G2458;
  assign new_G349 = ~new_G605;
  assign new_G350 = ~new_G608;
  assign new_G2265 = new_G2048 & new_G1998 & new_G1895 & new_G1947;
  assign new_G2273 = ~new_G1993 | ~new_G1895 | ~new_G1947;
  assign new_G2274 = ~new_G1895 | ~new_G1998 | ~new_G2043 | ~new_G1947;
  assign new_G2309 = new_G2262 & new_G2210 & new_G2103 & new_G2157;
  assign new_G2313 = ~new_G2205 | ~new_G2103 | ~new_G2157;
  assign new_G2314 = ~new_G2103 | ~new_G2210 | ~new_G2257 | ~new_G2157;
  assign new_G2325 = new_G1947;
  assign new_G2372 = new_G2157;
  assign new_G2523 = ~new_G2444;
  assign new_G2533 = ~new_G2454;
  assign new_G3121 = new_G2317;
  assign new_G3131 = new_G2317;
  assign new_G3155 = new_G2338;
  assign new_G3163 = new_G2338;
  assign new_G3171 = new_G2351;
  assign new_G3179 = new_G2351;
  assign new_G3187 = new_G2364;
  assign new_G3197 = new_G2364;
  assign new_G3221 = new_G2380;
  assign new_G3229 = new_G2380;
  assign new_G3237 = new_G2388;
  assign new_G3245 = new_G2388;
  assign G351 = ~new_G349 | ~new_G350;
  assign new_G2275 = ~new_G2274 | ~new_G2273 | ~new_G2271 | ~new_G2272;
  assign new_G2315 = ~new_G2314 | ~new_G2313 | ~new_G2311 | ~new_G2312;
  assign new_G3329 = ~new_G3323;
  assign G372 = new_G2309 & new_G2265;
  assign new_G2324 = ~new_G3131 | ~new_G3138;
  assign new_G2350 = ~new_G3163 | ~new_G3170;
  assign new_G2363 = ~new_G3179 | ~new_G3186;
  assign new_G2371 = ~new_G3197 | ~new_G3204;
  assign new_G2387 = ~new_G3229 | ~new_G3236;
  assign new_G2400 = ~new_G3245 | ~new_G3252;
  assign new_G2268 = new_G2265;
  assign new_G3137 = ~new_G3131;
  assign new_G3161 = ~new_G3155;
  assign new_G2345 = ~new_G3155 | ~new_G3162;
  assign new_G3169 = ~new_G3163;
  assign new_G3177 = ~new_G3171;
  assign new_G2358 = ~new_G3171 | ~new_G3178;
  assign new_G3185 = ~new_G3179;
  assign new_G3203 = ~new_G3197;
  assign new_G3235 = ~new_G3229;
  assign new_G3243 = ~new_G3237;
  assign new_G2395 = ~new_G3237 | ~new_G3244;
  assign new_G3251 = ~new_G3245;
  assign new_G3227 = ~new_G3221;
  assign new_G2432 = ~new_G3221 | ~new_G3228;
  assign new_G2490 = new_G2309 & new_G2485;
  assign new_G3127 = ~new_G3121;
  assign new_G3130 = ~new_G3121 | ~new_G3128;
  assign new_G3139 = new_G2325;
  assign new_G3147 = new_G2325;
  assign new_G3193 = ~new_G3187;
  assign new_G3196 = ~new_G3187 | ~new_G3194;
  assign new_G3205 = new_G2372;
  assign new_G3213 = new_G2372;
  assign new_G2307 = ~new_G2265 | ~new_G2315;
  assign new_G2308 = ~new_G2275;
  assign new_G2323 = ~new_G3134 | ~new_G3137;
  assign new_G2349 = ~new_G3166 | ~new_G3169;
  assign new_G2362 = ~new_G3182 | ~new_G3185;
  assign new_G2370 = ~new_G3200 | ~new_G3203;
  assign new_G2386 = ~new_G3232 | ~new_G3235;
  assign new_G2399 = ~new_G3248 | ~new_G3251;
  assign new_G2344 = ~new_G3158 | ~new_G3161;
  assign new_G2357 = ~new_G3174 | ~new_G3177;
  assign new_G2394 = ~new_G3240 | ~new_G3243;
  assign new_G2431 = ~new_G3224 | ~new_G3227;
  assign new_G2464 = new_G2315 & new_G2302;
  assign new_G2491 = new_G2489 | new_G2490;
  assign new_G3129 = ~new_G3124 | ~new_G3127;
  assign new_G3195 = ~new_G3190 | ~new_G3193;
  assign new_G368 = new_G2307 & new_G2308;
  assign new_G1615 = ~new_G2323 | ~new_G2324;
  assign new_G2337 = ~new_G3147 | ~new_G3154;
  assign new_G1633 = ~new_G2349 | ~new_G2350;
  assign new_G1642 = ~new_G2362 | ~new_G2363;
  assign new_G1651 = ~new_G2370 | ~new_G2371;
  assign new_G2379 = ~new_G3213 | ~new_G3220;
  assign new_G1669 = ~new_G2386 | ~new_G2387;
  assign new_G1678 = ~new_G2399 | ~new_G2400;
  assign new_G3145 = ~new_G3139;
  assign new_G2332 = ~new_G3139 | ~new_G3146;
  assign new_G3153 = ~new_G3147;
  assign new_G2346 = ~new_G2344 | ~new_G2345;
  assign new_G2359 = ~new_G2357 | ~new_G2358;
  assign new_G3219 = ~new_G3213;
  assign new_G2396 = ~new_G2394 | ~new_G2395;
  assign new_G3211 = ~new_G3205;
  assign new_G2425 = ~new_G3205 | ~new_G3212;
  assign new_G2433 = ~new_G2431 | ~new_G2432;
  assign new_G3272 = ~new_G3129 | ~new_G3130;
  assign new_G3308 = ~new_G3195 | ~new_G3196;
  assign G369 = ~new_G368;
  assign new_G1613 = ~new_G1615;
  assign new_G2336 = ~new_G3150 | ~new_G3153;
  assign new_G1631 = ~new_G1633;
  assign new_G1640 = ~new_G1642;
  assign new_G1649 = ~new_G1651;
  assign new_G2378 = ~new_G3216 | ~new_G3219;
  assign new_G1667 = ~new_G1669;
  assign new_G1676 = ~new_G1678;
  assign new_G2331 = ~new_G3142 | ~new_G3145;
  assign new_G2424 = ~new_G3208 | ~new_G3211;
  assign new_G2467 = new_G2464;
  assign new_G2495 = new_G2491;
  assign new_G3295 = new_G2464;
  assign new_G3374 = G330 & new_G2491;
  assign new_G1614 = new_G1613 & new_G1610;
  assign new_G1624 = ~new_G2336 | ~new_G2337;
  assign new_G1632 = new_G1631 & new_G1628;
  assign new_G1641 = new_G1640 & new_G1637;
  assign new_G1650 = new_G1649 & new_G1646;
  assign new_G1660 = ~new_G2378 | ~new_G2379;
  assign new_G1668 = new_G1667 & new_G1664;
  assign new_G1677 = new_G1676 & new_G1673;
  assign new_G2333 = ~new_G2331 | ~new_G2332;
  assign new_G2406 = new_G2346;
  assign new_G2409 = new_G2346;
  assign new_G2415 = new_G2359;
  assign new_G2419 = new_G2359;
  assign new_G2426 = ~new_G2424 | ~new_G2425;
  assign new_G2439 = new_G2396;
  assign new_G2518 = new_G2433 & new_G2461;
  assign new_G3276 = ~new_G3272;
  assign new_G3312 = ~new_G3308;
  assign new_G2612 = G330 & new_G2396;
  assign new_G3326 = new_G2433;
  assign new_G1617 = ~new_G1616 & ~new_G1612 & ~new_G1614;
  assign new_G1622 = ~new_G1624;
  assign new_G1635 = ~new_G1634 & ~new_G1630 & ~new_G1632;
  assign new_G1644 = ~new_G1643 & ~new_G1639 & ~new_G1641;
  assign new_G1653 = ~new_G1652 & ~new_G1648 & ~new_G1650;
  assign new_G1658 = ~new_G1660;
  assign new_G1671 = ~new_G1670 & ~new_G1666 & ~new_G1668;
  assign new_G1680 = ~new_G1679 & ~new_G1675 & ~new_G1677;
  assign new_G2500 = new_G2467 & new_G2268;
  assign new_G2505 = new_G2495 & new_G2268;
  assign new_G2519 = new_G2455 | new_G2518;
  assign new_G3378 = ~new_G3374;
  assign new_G2642 = ~new_G2467;
  assign new_G2645 = new_G2467;
  assign new_G3301 = ~new_G3295;
  assign new_G1623 = new_G1622 & new_G1619;
  assign new_G1659 = new_G1658 & new_G1655;
  assign new_G2401 = new_G2333;
  assign new_G2501 = new_G2275 | new_G2500;
  assign new_G2511 = new_G2409 & new_G2495 & new_G2419;
  assign new_G2512 = new_G2495 & new_G2415;
  assign new_G2513 = new_G2426 & new_G2439 & new_G2433;
  assign new_G2514 = new_G2439 & new_G2433;
  assign new_G2517 = new_G2467 & new_G2415;
  assign new_G2531 = ~new_G2409 | ~new_G2451;
  assign new_G2532 = ~new_G2467 | ~new_G2409 | ~new_G2419;
  assign new_G2534 = ~new_G2426 | ~new_G2455;
  assign new_G2535 = ~new_G2461 | ~new_G2426 | ~new_G2433;
  assign new_G2607 = ~new_G3326 | ~new_G3329;
  assign new_G3330 = ~new_G3326;
  assign new_G2643 = new_G2642 & G330 & new_G2491;
  assign new_G2687 = new_G1617 & new_G2680;
  assign new_G2725 = new_G1635 & new_G2718;
  assign new_G2742 = new_G1644 & new_G2735;
  assign new_G2760 = new_G1653 & new_G2753;
  assign new_G2794 = new_G1671 & new_G2787;
  assign new_G2811 = new_G1680 & new_G2804;
  assign new_G3280 = new_G2333;
  assign new_G3290 = new_G2409;
  assign new_G3298 = new_G2415;
  assign new_G3316 = new_G2426;
  assign new_G3406 = new_G2612;
  assign new_G3414 = new_G2612;
  assign new_G3422 = new_G2439 & new_G2439;
  assign new_G1626 = ~new_G1625 & ~new_G1621 & ~new_G1623;
  assign new_G1662 = ~new_G1661 & ~new_G1657 & ~new_G1659;
  assign new_G2567 = G330 & new_G2512;
  assign new_G2589 = G330 & new_G2513;
  assign new_G2608 = ~new_G3323 | ~new_G3330;
  assign new_G2654 = new_G2519;
  assign new_G3253 = new_G2505;
  assign new_G3277 = ~new_G2532 | ~new_G2530 | ~new_G2531;
  assign new_G3287 = new_G2448 | new_G2517;
  assign new_G3305 = ~new_G2535 | ~new_G2533 | ~new_G2534;
  assign new_G3313 = new_G2519;
  assign new_G3350 = G330 & new_G2511;
  assign new_G932 = new_G2643 | new_G2645;
  assign new_G2508 = new_G2419 & new_G2409 & new_G2495 & new_G2401;
  assign new_G2524 = ~new_G2401 | ~new_G2445;
  assign new_G2525 = ~new_G2451 | ~new_G2401 | ~new_G2406;
  assign new_G2526 = ~new_G2467 | ~new_G2419 | ~new_G2401 | ~new_G2406;
  assign new_G3294 = ~new_G3290;
  assign new_G2609 = ~new_G2607 | ~new_G2608;
  assign new_G3410 = ~new_G3406;
  assign new_G3418 = ~new_G3414;
  assign new_G2624 = ~new_G3422 | ~new_G3425;
  assign new_G3426 = ~new_G3422;
  assign new_G2629 = new_G2501;
  assign new_G2647 = ~new_G2643 & ~new_G2645;
  assign new_G2706 = new_G1626 & new_G2699;
  assign new_G2777 = new_G1662 & new_G2770;
  assign new_G3264 = new_G2501;
  assign new_G3284 = ~new_G3280;
  assign new_G3302 = ~new_G3298;
  assign new_G3303 = ~new_G3298 | ~new_G3301;
  assign new_G3320 = ~new_G3316;
  assign new_G3398 = G330 & new_G2514;
  assign new_G2657 = ~new_G2654;
  assign new_G398 = new_G2519 & new_G2654;
  assign new_G933 = new_G932 & new_G927;
  assign new_G2527 = ~new_G2526 | ~new_G2525 | ~new_G2523 | ~new_G2524;
  assign new_G3259 = ~new_G3253;
  assign new_G3354 = ~new_G3350;
  assign new_G3293 = ~new_G3287;
  assign new_G2563 = ~new_G3287 | ~new_G3294;
  assign new_G3311 = ~new_G3305;
  assign new_G2585 = ~new_G3305 | ~new_G3312;
  assign new_G2625 = ~new_G3419 | ~new_G3426;
  assign new_G3283 = ~new_G3277;
  assign new_G3286 = ~new_G3277 | ~new_G3284;
  assign new_G3304 = ~new_G3295 | ~new_G3302;
  assign new_G3319 = ~new_G3313;
  assign new_G3322 = ~new_G3313 | ~new_G3320;
  assign new_G3358 = new_G2567;
  assign new_G3366 = new_G2567;
  assign new_G3382 = new_G2589;
  assign new_G3390 = new_G2589;
  assign new_G397 = new_G2657 & G330 & new_G2514;
  assign new_G2544 = G330 & new_G2508;
  assign new_G2562 = ~new_G3290 | ~new_G3293;
  assign new_G2584 = ~new_G3308 | ~new_G3311;
  assign new_G3402 = ~new_G3398;
  assign new_G2626 = ~new_G2624 | ~new_G2625;
  assign new_G2632 = ~new_G2629;
  assign new_G2634 = new_G2501 & new_G2629;
  assign new_G2650 = new_G2647;
  assign new_G3268 = ~new_G3264;
  assign new_G3256 = new_G2508;
  assign new_G3285 = ~new_G3280 | ~new_G3283;
  assign new_G3321 = ~new_G3316 | ~new_G3319;
  assign new_G3371 = ~new_G3303 | ~new_G3304;
  assign new_G3403 = new_G2609;
  assign new_G3411 = new_G2609;
  assign new_G362 = new_G938 | new_G929 | new_G933;
  assign new_G1030 = ~new_G938 & ~new_G929 & ~new_G933;
  assign G399 = new_G397 | new_G398;
  assign new_G2564 = ~new_G2562 | ~new_G2563;
  assign new_G3362 = ~new_G3358;
  assign new_G3370 = ~new_G3366;
  assign new_G2586 = ~new_G2584 | ~new_G2585;
  assign new_G3386 = ~new_G3382;
  assign new_G3394 = ~new_G3390;
  assign new_G2633 = new_G2632 & G330 & new_G2505;
  assign new_G3261 = new_G2527;
  assign new_G3269 = new_G2527;
  assign new_G3347 = ~new_G3285 | ~new_G3286;
  assign new_G3395 = ~new_G3321 | ~new_G3322;
  assign new_G363 = ~new_G1030;
  assign new_G2536 = ~new_G3256 | ~new_G3259;
  assign new_G3260 = ~new_G3256;
  assign new_G3377 = ~new_G3371;
  assign new_G2580 = ~new_G3371 | ~new_G3378;
  assign new_G3409 = ~new_G3403;
  assign new_G2616 = ~new_G3403 | ~new_G3410;
  assign new_G3417 = ~new_G3411;
  assign new_G2622 = ~new_G3411 | ~new_G3418;
  assign new_G2635 = ~new_G2633 & ~new_G2634;
  assign new_G2805 = new_G2626 & new_G2802;
  assign new_G2808 = new_G2626 & new_G2803;
  assign new_G3334 = new_G2544;
  assign new_G3342 = new_G2544;
  assign new_G3454 = new_G2650;
  assign G364 = new_G362 & new_G363;
  assign new_G2537 = ~new_G3253 | ~new_G3260;
  assign new_G3275 = ~new_G3269;
  assign new_G2540 = ~new_G3269 | ~new_G3276;
  assign new_G3353 = ~new_G3347;
  assign new_G2557 = ~new_G3347 | ~new_G3354;
  assign new_G2579 = ~new_G3374 | ~new_G3377;
  assign new_G3401 = ~new_G3395;
  assign new_G2602 = ~new_G3395 | ~new_G3402;
  assign new_G2615 = ~new_G3406 | ~new_G3409;
  assign new_G2621 = ~new_G3414 | ~new_G3417;
  assign new_G3267 = ~new_G3261;
  assign new_G3112 = ~new_G3261 | ~new_G3268;
  assign new_G3355 = new_G2564;
  assign new_G3363 = new_G2564;
  assign new_G3379 = new_G2586;
  assign new_G3387 = new_G2586;
  assign new_G2538 = ~new_G2536 | ~new_G2537;
  assign new_G2539 = ~new_G3272 | ~new_G3275;
  assign new_G3338 = ~new_G3334;
  assign new_G3346 = ~new_G3342;
  assign new_G2556 = ~new_G3350 | ~new_G3353;
  assign new_G2581 = ~new_G2579 | ~new_G2580;
  assign new_G2601 = ~new_G3398 | ~new_G3401;
  assign new_G2617 = ~new_G2615 | ~new_G2616;
  assign new_G2623 = ~new_G2621 | ~new_G2622;
  assign new_G2638 = new_G2635;
  assign new_G3458 = ~new_G3454;
  assign new_G2814 = new_G2811 | new_G2805 | new_G2808;
  assign new_G2816 = ~new_G2811 & ~new_G2805 & ~new_G2808;
  assign new_G3111 = ~new_G3264 | ~new_G3267;
  assign new_G2541 = ~new_G2539 | ~new_G2540;
  assign new_G2558 = ~new_G2556 | ~new_G2557;
  assign new_G3361 = ~new_G3355;
  assign new_G2571 = ~new_G3355 | ~new_G3362;
  assign new_G3369 = ~new_G3363;
  assign new_G2577 = ~new_G3363 | ~new_G3370;
  assign new_G3385 = ~new_G3379;
  assign new_G2593 = ~new_G3379 | ~new_G3386;
  assign new_G3393 = ~new_G3387;
  assign new_G2598 = ~new_G3387 | ~new_G3394;
  assign new_G2603 = ~new_G2601 | ~new_G2602;
  assign new_G3113 = ~new_G3111 | ~new_G3112;
  assign new_G3116 = G330 & new_G2538;
  assign new_G3451 = ~new_G2623;
  assign new_G395 = ~new_G2816;
  assign new_G2570 = ~new_G3358 | ~new_G3361;
  assign new_G2576 = ~new_G3366 | ~new_G3369;
  assign new_G2592 = ~new_G3382 | ~new_G3385;
  assign new_G2597 = ~new_G3390 | ~new_G3393;
  assign new_G2736 = new_G2581 & new_G2733;
  assign new_G2739 = new_G2581 & new_G2734;
  assign new_G2788 = new_G2617 & new_G2785;
  assign new_G3438 = new_G2638;
  assign new_G3446 = new_G2617 & new_G2647;
  assign new_G3459 = new_G2814;
  assign G396 = new_G2814 & new_G395;
  assign new_G3119 = ~new_G3113;
  assign new_G3120 = ~new_G3116;
  assign new_G2572 = ~new_G2570 | ~new_G2571;
  assign new_G2578 = ~new_G2576 | ~new_G2577;
  assign new_G2594 = ~new_G2592 | ~new_G2593;
  assign new_G2599 = ~new_G2597 | ~new_G2598;
  assign new_G2677 = ~new_G3451 | ~new_G3458;
  assign new_G3457 = ~new_G3451;
  assign new_G2700 = new_G2558 & new_G2697;
  assign new_G2771 = new_G2603 & new_G2768;
  assign new_G3331 = new_G2541;
  assign new_G3339 = new_G2541;
  assign new_G3427 = new_G2558;
  assign new_G3443 = new_G2603;
  assign new_G954 = ~new_G3116 | ~new_G3119;
  assign new_G955 = ~new_G3113 | ~new_G3120;
  assign new_G2600 = ~new_G2599;
  assign new_G3442 = ~new_G3438;
  assign new_G3450 = ~new_G3446;
  assign new_G2676 = ~new_G3454 | ~new_G3457;
  assign new_G2745 = new_G2742 | new_G2736 | new_G2739;
  assign new_G2748 = ~new_G2742 & ~new_G2736 & ~new_G2739;
  assign new_G3465 = ~new_G3459;
  assign new_G3435 = ~new_G2578;
  assign new_G950 = ~new_G954 | ~new_G955;
  assign new_G3337 = ~new_G3331;
  assign new_G2548 = ~new_G3331 | ~new_G3338;
  assign new_G3345 = ~new_G3339;
  assign new_G2553 = ~new_G3339 | ~new_G3346;
  assign new_G2661 = ~new_G2600 & ~new_G2650;
  assign new_G2662 = new_G2650 & new_G2594 & new_G2617 & new_G2603;
  assign new_G3433 = ~new_G3427;
  assign new_G3449 = ~new_G3443;
  assign new_G2672 = ~new_G3443 | ~new_G3450;
  assign new_G2674 = ~new_G2676 | ~new_G2677;
  assign new_G2719 = new_G2572 & new_G2716;
  assign new_G2754 = new_G2594 & new_G2751;
  assign new_G3430 = new_G2572 & new_G2635;
  assign new_G383 = ~new_G2748;
  assign new_G951 = new_G950 & new_G943;
  assign new_G2547 = ~new_G3334 | ~new_G3337;
  assign new_G2552 = ~new_G3342 | ~new_G3345;
  assign new_G2663 = new_G2661 | new_G2662;
  assign new_G2670 = ~new_G3435 | ~new_G3442;
  assign new_G3441 = ~new_G3435;
  assign new_G2671 = ~new_G3446 | ~new_G3449;
  assign new_G2675 = ~new_G2674;
  assign new_G3491 = new_G2745;
  assign new_G3499 = new_G2745;
  assign G384 = new_G2745 & new_G383;
  assign new_G2549 = ~new_G2547 | ~new_G2548;
  assign new_G2554 = ~new_G2552 | ~new_G2553;
  assign new_G2664 = ~new_G3430 | ~new_G3433;
  assign new_G3434 = ~new_G3430;
  assign new_G2669 = ~new_G3438 | ~new_G3441;
  assign new_G2673 = ~new_G2671 | ~new_G2672;
  assign new_G2757 = new_G2663 & new_G2752;
  assign new_G2791 = new_G2675 & new_G2786;
  assign new_G365 = new_G951 | new_G944 | new_G947;
  assign new_G1031 = ~new_G951 & ~new_G944 & ~new_G947;
  assign new_G2555 = ~new_G2554;
  assign new_G2665 = ~new_G3427 | ~new_G3434;
  assign new_G2667 = ~new_G2669 | ~new_G2670;
  assign new_G2774 = new_G2673 & new_G2769;
  assign new_G3497 = ~new_G3491;
  assign new_G3505 = ~new_G3499;
  assign new_G366 = ~new_G1031;
  assign new_G2658 = ~new_G2555 & ~new_G2638;
  assign new_G2659 = new_G2638 & new_G2549 & new_G2572 & new_G2558;
  assign new_G2666 = ~new_G2664 | ~new_G2665;
  assign new_G2668 = ~new_G2667;
  assign new_G2681 = new_G2549 & new_G2678;
  assign new_G2763 = new_G2760 | new_G2754 | new_G2757;
  assign new_G2765 = ~new_G2760 & ~new_G2754 & ~new_G2757;
  assign new_G2797 = new_G2794 | new_G2788 | new_G2791;
  assign new_G2799 = ~new_G2794 & ~new_G2788 & ~new_G2791;
  assign G367 = new_G365 & new_G366;
  assign new_G2660 = new_G2658 | new_G2659;
  assign new_G2703 = new_G2666 & new_G2698;
  assign new_G2722 = new_G2668 & new_G2717;
  assign new_G2780 = new_G2777 | new_G2771 | new_G2774;
  assign new_G2782 = ~new_G2777 & ~new_G2771 & ~new_G2774;
  assign new_G386 = ~new_G2765;
  assign new_G392 = ~new_G2799;
  assign new_G2684 = new_G2660 & new_G2679;
  assign new_G3462 = new_G2797;
  assign new_G3470 = new_G2763;
  assign G387 = new_G2763 & new_G386;
  assign new_G389 = ~new_G2782;
  assign G393 = new_G2797 & new_G392;
  assign new_G2709 = new_G2706 | new_G2700 | new_G2703;
  assign new_G2713 = ~new_G2706 & ~new_G2700 & ~new_G2703;
  assign new_G2728 = new_G2725 | new_G2719 | new_G2722;
  assign new_G2730 = ~new_G2725 & ~new_G2719 & ~new_G2722;
  assign new_G2922 = new_G2765 & new_G2782 & new_G2816 & new_G2799;
  assign new_G3467 = new_G2780;
  assign G390 = new_G2780 & new_G389;
  assign new_G2690 = new_G2687 | new_G2681 | new_G2684;
  assign new_G2694 = ~new_G2687 & ~new_G2681 & ~new_G2684;
  assign new_G2821 = ~new_G3462 | ~new_G3465;
  assign new_G3466 = ~new_G3462;
  assign new_G3474 = ~new_G3470;
  assign G378 = new_G2709 & new_G2709;
  assign new_G380 = ~new_G2730;
  assign new_G2822 = ~new_G3459 | ~new_G3466;
  assign new_G3473 = ~new_G3467;
  assign new_G2827 = ~new_G3467 | ~new_G3474;
  assign new_G2839 = new_G2728;
  assign new_G2883 = new_G2709 & new_G2871;
  assign new_G3507 = new_G2709;
  assign G375 = new_G2690 & new_G2690;
  assign G381 = new_G2728 & new_G380;
  assign new_G2823 = ~new_G2821 | ~new_G2822;
  assign new_G2826 = ~new_G3470 | ~new_G3473;
  assign new_G2880 = new_G2871 & new_G2690;
  assign new_G2925 = new_G2694 & new_G2713 & new_G2748 & new_G2730;
  assign new_G2928 = new_G2874 & new_G2713 & new_G2694;
  assign new_G3510 = new_G2690;
  assign new_G2828 = ~new_G2826 | ~new_G2827;
  assign new_G3494 = new_G2839;
  assign new_G3502 = new_G2839;
  assign new_G3513 = ~new_G3507;
  assign new_G3544 = new_G2883;
  assign new_G3552 = new_G2883;
  assign new_G406 = new_G2922 & new_G2925;
  assign new_G2929 = new_G2922 & new_G2925;
  assign new_G3475 = new_G2823;
  assign new_G3483 = new_G2823;
  assign new_G3514 = ~new_G3510;
  assign new_G3515 = ~new_G3510 | ~new_G3513;
  assign new_G3541 = new_G2880;
  assign new_G3549 = new_G2880;
  assign G407 = ~new_G406;
  assign new_G2930 = ~new_G2928 & ~new_G2929;
  assign new_G2842 = ~new_G3494 | ~new_G3497;
  assign new_G3498 = ~new_G3494;
  assign new_G2852 = ~new_G3502 | ~new_G3505;
  assign new_G3506 = ~new_G3502;
  assign new_G3548 = ~new_G3544;
  assign new_G3556 = ~new_G3552;
  assign new_G3478 = new_G2828;
  assign new_G3486 = new_G2828;
  assign new_G3516 = ~new_G3507 | ~new_G3514;
  assign new_G408 = G213 & new_G2930;
  assign new_G3481 = ~new_G3475;
  assign new_G3489 = ~new_G3483;
  assign new_G2843 = ~new_G3491 | ~new_G3498;
  assign new_G2853 = ~new_G3499 | ~new_G3506;
  assign new_G3547 = ~new_G3541;
  assign new_G2887 = ~new_G3541 | ~new_G3548;
  assign new_G2896 = ~new_G3549 | ~new_G3556;
  assign new_G3555 = ~new_G3549;
  assign new_G3520 = ~new_G3515 | ~new_G3516;
  assign G409 = ~new_G408;
  assign new_G2831 = ~new_G3478 | ~new_G3481;
  assign new_G3482 = ~new_G3478;
  assign new_G2836 = ~new_G3486 | ~new_G3489;
  assign new_G3490 = ~new_G3486;
  assign new_G2844 = ~new_G2842 | ~new_G2843;
  assign new_G2848 = ~new_G2852 | ~new_G2853;
  assign new_G2886 = ~new_G3544 | ~new_G3547;
  assign new_G2895 = ~new_G3552 | ~new_G3555;
  assign new_G2832 = ~new_G3475 | ~new_G3482;
  assign new_G2837 = ~new_G3483 | ~new_G3490;
  assign new_G2849 = ~new_G2848;
  assign new_G3524 = ~new_G3520;
  assign new_G2888 = ~new_G2886 | ~new_G2887;
  assign new_G2891 = ~new_G2895 | ~new_G2896;
  assign new_G2833 = ~new_G2831 | ~new_G2832;
  assign new_G2838 = ~new_G2836 | ~new_G2837;
  assign new_G2892 = ~new_G2891;
  assign new_G3517 = new_G2844;
  assign new_G2906 = new_G2900 & new_G2844 & new_G2888;
  assign new_G2908 = new_G2903 & new_G2849 & new_G2888;
  assign new_G2913 = ~new_G2838;
  assign new_G3523 = ~new_G3517;
  assign new_G2855 = ~new_G3517 | ~new_G3524;
  assign new_G2907 = new_G2903 & new_G2844 & new_G2892;
  assign new_G2909 = new_G2900 & new_G2849 & new_G2892;
  assign new_G3525 = new_G2833;
  assign new_G3533 = new_G2833;
  assign new_G2854 = ~new_G3520 | ~new_G3523;
  assign new_G2910 = new_G2909 | new_G2908 | new_G2906 | new_G2907;
  assign new_G3560 = new_G2913;
  assign new_G3568 = new_G2913;
  assign new_G2856 = ~new_G2854 | ~new_G2855;
  assign new_G3539 = ~new_G3533;
  assign new_G3531 = ~new_G3525;
  assign new_G3572 = ~new_G3568;
  assign new_G3564 = ~new_G3560;
  assign new_G3557 = new_G2910;
  assign new_G3565 = new_G2910;
  assign new_G3528 = new_G2856;
  assign new_G3536 = new_G2856;
  assign new_G2921 = ~new_G3557 | ~new_G3564;
  assign new_G2917 = ~new_G3565 | ~new_G3572;
  assign new_G3571 = ~new_G3565;
  assign new_G3563 = ~new_G3557;
  assign new_G2863 = ~new_G3528 | ~new_G3531;
  assign new_G2859 = ~new_G3536 | ~new_G3539;
  assign new_G2920 = ~new_G3560 | ~new_G3563;
  assign new_G2916 = ~new_G3568 | ~new_G3571;
  assign new_G3540 = ~new_G3536;
  assign new_G3532 = ~new_G3528;
  assign new_G2864 = ~new_G3525 | ~new_G3532;
  assign new_G2860 = ~new_G3533 | ~new_G3540;
  assign new_G403 = ~new_G2920 | ~new_G2921;
  assign new_G404 = ~new_G2916 | ~new_G2917;
  assign new_G400 = ~new_G2863 | ~new_G2864;
  assign new_G401 = ~new_G2859 | ~new_G2860;
  assign G405 = new_G403 & new_G404;
  assign G402 = ~new_G400 | ~new_G401;
endmodule
