// Benchmark "./benchmarks/iscas85/c7552" written by ABC on Sun Apr 28 12:32:39 2024

module c7552  ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496,
    G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253,
    G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743,
    G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432,
    G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_G400, new_G1184, new_G1501, new_G2857, new_G4442, new_G4514,
    new_G401, new_G573, new_G574, new_G575, new_G1178, new_G1186,
    new_G1192, new_G1198, new_G1205, new_G1206, new_G1207, new_G1210,
    new_G1458, new_G1461, new_G1464, new_G1471, new_G1475, new_G1482,
    new_G1488, new_G1495, new_G1499, new_G1500, new_G1503, new_G1512,
    new_G1518, new_G1524, new_G1535, new_G1541, new_G2207, new_G2210,
    new_G2213, new_G2220, new_G2226, new_G2232, new_G2238, new_G2241,
    new_G2249, new_G2255, new_G2258, new_G2828, new_G3700, new_G3703,
    new_G3707, new_G3713, new_G3719, new_G3725, new_G3731, new_G3739,
    new_G3745, new_G3751, new_G4121, new_G4396, new_G4402, new_G4407,
    new_G4412, new_G4417, new_G4422, new_G4429, new_G4434, new_G4439,
    new_G4833, new_G2876, new_G2878, new_G1519, new_G2871, new_G2883,
    new_G280, new_G4839, new_G572, new_G581, new_G587, new_G601, new_G606,
    new_G650, new_G657, new_G671, new_G678, new_G777, new_G1115, new_G1336,
    new_G1350, new_G1477, new_G1507, new_G1514, new_G1530, new_G2259,
    new_G2833, new_G2872, new_G2886, new_G2892, new_G2905, new_G2909,
    new_G3622, new_G3635, new_G3755, new_G4640, new_G4653, new_G4873,
    new_G4876, new_G4881, new_G4889, new_G4905, new_G4916, new_G4921,
    new_G5175, new_G5178, new_G5186, new_G5191, new_G5199, new_G5215,
    new_G5223, new_G5393, new_G5401, new_G5409, new_G5417, new_G5425,
    new_G5433, new_G5441, new_G5449, new_G5457, new_G5745, new_G5753,
    new_G5761, new_G5769, new_G5777, new_G5785, new_G5793, new_G5801,
    new_G5809, new_G5865, new_G5873, new_G5881, new_G5889, new_G5897,
    new_G5905, new_G5913, new_G5921, new_G5985, new_G5993, new_G6001,
    new_G6009, new_G6017, new_G6025, new_G6033, new_G6041, new_G6514,
    new_G6554, new_G6567, new_G6575, new_G6583, new_G6591, new_G6599,
    new_G6607, new_G6615, new_G6623, new_G6631, new_G6853, new_G6861,
    new_G6869, new_G6877, new_G6885, new_G6893, new_G6901, new_G6909,
    new_G6917, new_G784, new_G1014, new_G3221, new_G4913, new_G4929,
    new_G5183, new_G5231, new_G6511, new_G615, new_G594, new_G611,
    new_G617, new_G619, new_G621, new_G623, new_G625, new_G627, new_G664,
    new_G685, new_G691, new_G693, new_G695, new_G697, new_G699, new_G701,
    new_G703, new_G705, new_G707, new_G709, new_G4879, new_G4880,
    new_G4887, new_G4895, new_G4911, new_G4920, new_G4927, new_G5181,
    new_G5182, new_G5190, new_G5197, new_G5205, new_G5221, new_G5229,
    new_G1343, new_G1357, new_G1364, new_G1366, new_G1368, new_G1370,
    new_G1372, new_G1374, new_G1376, new_G1378, new_G1380, new_G1382,
    new_G5399, new_G5407, new_G5415, new_G5423, new_G5431, new_G5439,
    new_G5447, new_G5455, new_G5463, new_G5751, new_G5759, new_G5767,
    new_G5775, new_G5783, new_G5791, new_G5799, new_G5807, new_G5815,
    new_G2019, new_G2032, new_G2117, new_G2130, new_G2266, new_G2272,
    new_G2286, new_G2288, new_G2290, new_G2292, new_G2294, new_G5871,
    new_G5879, new_G5887, new_G5895, new_G5903, new_G5911, new_G5919,
    new_G5927, new_G5991, new_G5999, new_G6007, new_G6015, new_G6023,
    new_G6031, new_G6039, new_G6047, new_G2899, new_G2914, new_G2919,
    new_G2921, new_G2923, new_G2925, new_G2927, new_G2929, new_G2931,
    new_G6518, new_G3173, new_G6558, new_G6573, new_G6581, new_G6589,
    new_G6597, new_G6605, new_G6613, new_G6621, new_G6629, new_G6637,
    new_G3629, new_G3642, new_G3649, new_G3651, new_G3653, new_G3655,
    new_G3657, new_G3659, new_G3661, new_G3663, new_G3762, new_G3768,
    new_G3782, new_G3784, new_G3786, new_G3788, new_G3790, new_G6859,
    new_G6867, new_G6875, new_G6883, new_G6891, new_G6899, new_G6907,
    new_G6915, new_G6923, new_G4094, new_G4107, new_G4444, new_G4457,
    new_G4647, new_G4660, new_G4667, new_G4669, new_G4671, new_G4673,
    new_G4675, new_G4677, new_G4679, new_G4681, new_G4683, new_G4685,
    new_G4897, new_G5207, new_G6551, new_G763, new_G764, new_G4919,
    new_G886, new_G1005, new_G1006, new_G5189, new_G1018, new_G5237,
    new_G6517, new_G3169, new_G4935, new_G4970, new_G5239, new_G577,
    new_G616, new_G618, new_G620, new_G622, new_G624, new_G626, new_G628,
    new_G692, new_G694, new_G696, new_G698, new_G700, new_G702, new_G704,
    new_G706, new_G708, new_G710, new_G765, new_G4903, new_G885, new_G1007,
    new_G1017, new_G5213, new_G1363, new_G1365, new_G1367, new_G1369,
    new_G1371, new_G1373, new_G1375, new_G1377, new_G1379, new_G1381,
    new_G2026, new_G2039, new_G2046, new_G2048, new_G2050, new_G2052,
    new_G2054, new_G2056, new_G2058, new_G2060, new_G2062, new_G2064,
    new_G2124, new_G2137, new_G2144, new_G2146, new_G2148, new_G2150,
    new_G2152, new_G2154, new_G2156, new_G2158, new_G2160, new_G2162,
    new_G2279, new_G2285, new_G2287, new_G2289, new_G2291, new_G2293,
    new_G2296, new_G2298, new_G2300, new_G2302, new_G2304, new_G2918,
    new_G2920, new_G2922, new_G2924, new_G2926, new_G2928, new_G2930,
    new_G2932, new_G3168, new_G6557, new_G3211, new_G3648, new_G3650,
    new_G3652, new_G3654, new_G3656, new_G3658, new_G3660, new_G3662,
    new_G3665, new_G3666, new_G3775, new_G3781, new_G3783, new_G3785,
    new_G3787, new_G3789, new_G3792, new_G3794, new_G3796, new_G3798,
    new_G3800, new_G4101, new_G4114, new_G4123, new_G4126, new_G4129,
    new_G4132, new_G4135, new_G4138, new_G4141, new_G4144, new_G4147,
    new_G4150, new_G4451, new_G4464, new_G4471, new_G4473, new_G4475,
    new_G4477, new_G4479, new_G4481, new_G4483, new_G4485, new_G4487,
    new_G4489, new_G4666, new_G4668, new_G4670, new_G4672, new_G4674,
    new_G4676, new_G4678, new_G4680, new_G4682, new_G4684, new_G579,
    new_G629, new_G633, new_G637, new_G641, new_G645, new_G711, new_G715,
    new_G719, new_G723, new_G727, new_G731, new_G737, new_G745, new_G751,
    new_G757, new_G887, new_G1019, new_G5245, new_G1383, new_G1387,
    new_G1391, new_G1395, new_G1399, new_G1406, new_G1412, new_G1418,
    new_G2305, new_G2308, new_G2312, new_G2316, new_G2933, new_G2938,
    new_G2942, new_G2946, new_G2950, new_G3170, new_G3210, new_G3667,
    new_G3670, new_G3673, new_G3676, new_G3679, new_G3682, new_G3686,
    new_G3801, new_G3804, new_G3807, new_G3810, new_G3813, new_G4525,
    new_G4686, new_G4689, new_G4692, new_G4695, new_G4698, new_G4701,
    new_G4704, new_G4707, new_G4710, new_G4976, new_G5271, new_G5274,
    new_G5305, new_G5308, new_G5318, new_G6690, new_G6711, new_G6714,
    new_G7252, new_G7296, new_G7466, new_G907, new_G913, new_G915,
    new_G916, new_G1116, new_G2045, new_G2047, new_G2049, new_G2051,
    new_G2053, new_G2055, new_G2057, new_G2059, new_G2061, new_G2063,
    new_G2143, new_G2145, new_G2147, new_G2149, new_G2151, new_G2153,
    new_G2155, new_G2157, new_G2159, new_G2161, new_G2295, new_G2297,
    new_G2299, new_G2301, new_G2303, new_G3212, new_G3791, new_G3793,
    new_G3795, new_G3797, new_G3799, new_G4122, new_G4125, new_G4128,
    new_G4131, new_G4134, new_G4137, new_G4140, new_G4143, new_G4146,
    new_G4149, new_G4470, new_G4472, new_G4474, new_G4476, new_G4478,
    new_G4480, new_G4482, new_G4484, new_G4486, new_G4488, new_G4962,
    new_G5003, new_G5234, new_G5242, new_G5250, new_G5284, new_G802,
    new_G821, new_G845, new_G868, new_G877, new_G902, new_G908, new_G914,
    new_G917, new_G953, new_G1023, new_G1035, new_G1050, new_G1068,
    new_G1086, new_G1102, new_G1108, new_G1117, new_G5322, new_G1553,
    new_G1567, new_G1584, new_G1590, new_G1606, new_G1624, new_G1647,
    new_G1669, new_G1677, new_G1802, new_G1816, new_G1834, new_G1841,
    new_G1866, new_G1880, new_G1897, new_G1914, new_G1929, new_G2065,
    new_G2069, new_G2073, new_G2077, new_G2081, new_G2085, new_G2091,
    new_G2099, new_G2105, new_G2111, new_G2163, new_G2167, new_G2171,
    new_G2175, new_G2179, new_G2186, new_G2192, new_G2198, new_G2320,
    new_G2323, new_G2329, new_G2335, new_G2962, new_G2970, new_G2977,
    new_G2979, new_G2989, new_G2998, new_G3006, new_G3013, new_G3015,
    new_G3183, new_G3192, new_G3200, new_G3207, new_G3209, new_G3216,
    new_G3222, new_G6694, new_G3695, new_G3816, new_G3821, new_G3828,
    new_G3833, new_G3838, new_G4151, new_G4154, new_G4157, new_G4160,
    new_G4163, new_G4166, new_G4169, new_G4172, new_G4175, new_G7256,
    new_G7300, new_G4490, new_G4493, new_G4496, new_G4499, new_G4502,
    new_G4505, new_G4508, new_G4511, new_G7470, new_G4884, new_G4892,
    new_G4900, new_G4908, new_G4924, new_G4952, new_G4983, new_G4993,
    new_G5011, new_G5194, new_G5202, new_G5210, new_G5218, new_G5226,
    new_G5247, new_G5255, new_G5258, new_G5263, new_G5266, new_G5277,
    new_G5278, new_G5281, new_G5289, new_G5292, new_G5297, new_G5300,
    new_G5311, new_G5312, new_G5315, new_G5323, new_G5326, new_G5331,
    new_G5334, new_G5339, new_G5342, new_G5349, new_G5352, new_G5396,
    new_G5404, new_G5412, new_G5420, new_G5428, new_G5436, new_G5444,
    new_G5452, new_G5460, new_G5465, new_G5581, new_G5748, new_G5756,
    new_G5764, new_G5772, new_G5780, new_G5788, new_G5796, new_G5804,
    new_G5812, new_G5849, new_G5929, new_G6049, new_G6367, new_G6370,
    new_G6375, new_G6378, new_G6383, new_G6386, new_G6391, new_G6394,
    new_G6399, new_G6402, new_G6407, new_G6410, new_G6415, new_G6418,
    new_G6423, new_G6426, new_G6431, new_G6434, new_G6442, new_G6450,
    new_G6458, new_G6466, new_G6498, new_G6519, new_G6522, new_G6527,
    new_G6530, new_G6535, new_G6538, new_G6543, new_G6546, new_G6559,
    new_G6562, new_G6687, new_G6695, new_G6698, new_G6703, new_G6706,
    new_G6717, new_G6718, new_G6724, new_G6768, new_G7208, new_G7221,
    new_G7229, new_G7232, new_G7239, new_G7242, new_G7249, new_G7257,
    new_G7260, new_G7268, new_G7293, new_G7301, new_G7304, new_G7309,
    new_G7312, new_G7317, new_G7320, new_G7327, new_G7330, new_G7396,
    new_G7404, new_G7412, new_G7425, new_G7463, new_G7471, new_G7474,
    new_G7479, new_G7482, new_G7487, new_G7490, new_G7497, new_G7500,
    new_G7507, new_G7510, new_G7554, new_G1152, new_G5238, new_G1156,
    new_G5246, new_G5254, new_G5288, new_G3223, new_G4942, new_G4966,
    new_G5007, new_G5279, new_G5280, new_G5313, new_G5314, new_G6719,
    new_G6720, new_G790, new_G4888, new_G803, new_G4896, new_G825,
    new_G4904, new_G851, new_G4912, new_G893, new_G4928, new_G906,
    new_G912, new_G1024, new_G5198, new_G1036, new_G5206, new_G1053,
    new_G5214, new_G1072, new_G5222, new_G1091, new_G5230, new_G1112,
    new_G1121, new_G1153, new_G1157, new_G5253, new_G1216, new_G5261,
    new_G5262, new_G5269, new_G5270, new_G5287, new_G1239, new_G5295,
    new_G5296, new_G5303, new_G5304, new_G5321, new_G1262, new_G5329,
    new_G5330, new_G5337, new_G5338, new_G1544, new_G5400, new_G1554,
    new_G5408, new_G1571, new_G5416, new_G1596, new_G5424, new_G1607,
    new_G5432, new_G1628, new_G5440, new_G1653, new_G5448, new_G1685,
    new_G5456, new_G1693, new_G5464, new_G1793, new_G5752, new_G1803,
    new_G5760, new_G1820, new_G5768, new_G1848, new_G5776, new_G1857,
    new_G5784, new_G1867, new_G5792, new_G1883, new_G5800, new_G1901,
    new_G5808, new_G1919, new_G5816, new_G5855, new_G2351, new_G2366,
    new_G2384, new_G2391, new_G2417, new_G2431, new_G2448, new_G2465,
    new_G5935, new_G2597, new_G2612, new_G2629, new_G2635, new_G2652,
    new_G2670, new_G2693, new_G2715, new_G6055, new_G6373, new_G6374,
    new_G6381, new_G6382, new_G6389, new_G6390, new_G6397, new_G6398,
    new_G6405, new_G6406, new_G6413, new_G6414, new_G6421, new_G6422,
    new_G6429, new_G6430, new_G6437, new_G6438, new_G6446, new_G3059,
    new_G6454, new_G3068, new_G6462, new_G3076, new_G3079, new_G6470,
    new_G3090, new_G3099, new_G3107, new_G3114, new_G3116, new_G6502,
    new_G6525, new_G6526, new_G6533, new_G6534, new_G6541, new_G6542,
    new_G6549, new_G6550, new_G6565, new_G6566, new_G3220, new_G3292,
    new_G3308, new_G3327, new_G3335, new_G3362, new_G3376, new_G3393,
    new_G3410, new_G3425, new_G6693, new_G3503, new_G6701, new_G6702,
    new_G6709, new_G6710, new_G6728, new_G6772, new_G3853, new_G3868,
    new_G3885, new_G3891, new_G3908, new_G3926, new_G3949, new_G3971,
    new_G3979, new_G7212, new_G7227, new_G7255, new_G4202, new_G7263,
    new_G7264, new_G7272, new_G7299, new_G4225, new_G7307, new_G7308,
    new_G7315, new_G7316, new_G4297, new_G4305, new_G4312, new_G4314,
    new_G4324, new_G7400, new_G4333, new_G7408, new_G4341, new_G7416,
    new_G4348, new_G4349, new_G7431, new_G4389, new_G7469, new_G4530,
    new_G7477, new_G7478, new_G7485, new_G7486, new_G7513, new_G7514,
    new_G7558, new_G4932, new_G4956, new_G4973, new_G4987, new_G4997,
    new_G5017, new_G5099, new_G5345, new_G5346, new_G5355, new_G5356,
    new_G5372, new_G5380, new_G5471, new_G5523, new_G5587, new_G5669,
    new_G5857, new_G5868, new_G5876, new_G5884, new_G5892, new_G5900,
    new_G5908, new_G5916, new_G5924, new_G5969, new_G5988, new_G5996,
    new_G6004, new_G6012, new_G6020, new_G6028, new_G6036, new_G6044,
    new_G6057, new_G6439, new_G6447, new_G6455, new_G6463, new_G6471,
    new_G6474, new_G6479, new_G6482, new_G6487, new_G6490, new_G6495,
    new_G6503, new_G6506, new_G6570, new_G6578, new_G6586, new_G6594,
    new_G6602, new_G6610, new_G6618, new_G6626, new_G6634, new_G6671,
    new_G6721, new_G6729, new_G6732, new_G6737, new_G6740, new_G6745,
    new_G6748, new_G6755, new_G6758, new_G6765, new_G6773, new_G6776,
    new_G6781, new_G6784, new_G6789, new_G6792, new_G6799, new_G6802,
    new_G6832, new_G6856, new_G6864, new_G6872, new_G6880, new_G6888,
    new_G6896, new_G6904, new_G6912, new_G6920, new_G6925, new_G7041,
    new_G7205, new_G7213, new_G7216, new_G7224, new_G7235, new_G7236,
    new_G7245, new_G7246, new_G7265, new_G7273, new_G7276, new_G7283,
    new_G7286, new_G7323, new_G7324, new_G7333, new_G7334, new_G7361,
    new_G7364, new_G7369, new_G7372, new_G7377, new_G7380, new_G7385,
    new_G7388, new_G7393, new_G7401, new_G7409, new_G7417, new_G7420,
    new_G7428, new_G7493, new_G7494, new_G7503, new_G7504, new_G7515,
    new_G7518, new_G7523, new_G7526, new_G7531, new_G7534, new_G7541,
    new_G7544, new_G7551, new_G7559, new_G7562, new_G7567, new_G7570,
    new_G7575, new_G7578, new_G7585, new_G7588, new_G1176, new_G957,
    new_G791, new_G804, new_G826, new_G852, new_G894, new_G1025, new_G1037,
    new_G1054, new_G1073, new_G1092, new_G1154, new_G1158, new_G1215,
    new_G1224, new_G1225, new_G1233, new_G1234, new_G1238, new_G1247,
    new_G1248, new_G1256, new_G1257, new_G1261, new_G1270, new_G1271,
    new_G1279, new_G1280, new_G1545, new_G1555, new_G1572, new_G1597,
    new_G1608, new_G1629, new_G1654, new_G1686, new_G1694, new_G1794,
    new_G1804, new_G1821, new_G1849, new_G1858, new_G1868, new_G1884,
    new_G1902, new_G1920, new_G2954, new_G2955, new_G2963, new_G2964,
    new_G2971, new_G2972, new_G2980, new_G2981, new_G2990, new_G2991,
    new_G2999, new_G3000, new_G3007, new_G3008, new_G3016, new_G3017,
    new_G3019, new_G3020, new_G3174, new_G3175, new_G3184, new_G3185,
    new_G3193, new_G3194, new_G3201, new_G3202, new_G3213, new_G3214,
    new_G3227, new_G3502, new_G3511, new_G3512, new_G3520, new_G3521,
    new_G4201, new_G4210, new_G4211, new_G4224, new_G4233, new_G4234,
    new_G4242, new_G4243, new_G4529, new_G4538, new_G4539, new_G4547,
    new_G4548, new_G4552, new_G4553, new_G4946, new_G5347, new_G5348,
    new_G5357, new_G5358, new_G7237, new_G7238, new_G7247, new_G7248,
    new_G7325, new_G7326, new_G7335, new_G7336, new_G7495, new_G7496,
    new_G7505, new_G7506, new_G3244, new_G792, new_G805, new_G827,
    new_G853, new_G895, new_G1026, new_G1038, new_G1055, new_G1074,
    new_G1093, new_G1155, new_G1217, new_G1226, new_G1235, new_G1240,
    new_G1249, new_G1258, new_G1263, new_G1272, new_G1281, new_G5376,
    new_G5384, new_G1546, new_G1556, new_G1573, new_G1598, new_G1609,
    new_G1630, new_G1655, new_G1687, new_G1695, new_G1795, new_G1805,
    new_G1822, new_G1850, new_G1859, new_G1869, new_G1885, new_G1903,
    new_G1921, new_G5863, new_G2341, new_G5872, new_G2352, new_G5880,
    new_G2370, new_G5888, new_G2398, new_G5896, new_G2407, new_G5904,
    new_G2418, new_G5912, new_G2434, new_G5920, new_G2452, new_G5928,
    new_G2481, new_G5975, new_G2587, new_G5992, new_G2598, new_G6000,
    new_G2616, new_G6008, new_G2641, new_G6016, new_G2653, new_G6024,
    new_G2674, new_G6032, new_G2699, new_G6040, new_G2724, new_G2732,
    new_G6048, new_G2956, new_G2965, new_G2973, new_G2982, new_G2992,
    new_G3001, new_G3009, new_G3018, new_G3021, new_G6445, new_G3051,
    new_G6453, new_G3061, new_G6461, new_G3070, new_G6469, new_G3081,
    new_G6477, new_G6478, new_G6485, new_G6486, new_G6493, new_G6494,
    new_G6501, new_G3118, new_G6509, new_G6510, new_G3176, new_G3186,
    new_G3195, new_G3203, new_G3215, new_G3281, new_G6574, new_G3293,
    new_G6582, new_G3312, new_G6590, new_G3342, new_G6598, new_G3351,
    new_G6606, new_G3363, new_G6614, new_G3379, new_G6622, new_G3397,
    new_G6630, new_G3415, new_G6638, new_G6677, new_G3504, new_G3513,
    new_G3522, new_G6727, new_G3526, new_G6735, new_G6736, new_G6743,
    new_G6744, new_G6771, new_G3549, new_G6779, new_G6780, new_G6787,
    new_G6788, new_G6836, new_G3843, new_G6860, new_G3854, new_G6868,
    new_G3872, new_G6876, new_G3897, new_G6884, new_G3909, new_G6892,
    new_G3930, new_G6900, new_G3955, new_G6908, new_G3987, new_G6916,
    new_G3995, new_G6924, new_G7211, new_G4179, new_G7219, new_G7220,
    new_G4196, new_G7228, new_G4203, new_G4212, new_G7271, new_G4220,
    new_G4226, new_G4235, new_G4244, new_G7367, new_G7368, new_G7375,
    new_G7376, new_G7383, new_G7384, new_G7391, new_G7392, new_G7399,
    new_G4326, new_G7407, new_G4335, new_G7415, new_G4343, new_G7423,
    new_G7424, new_G4353, new_G7432, new_G4531, new_G4540, new_G4549,
    new_G4554, new_G7521, new_G7522, new_G7529, new_G7530, new_G7557,
    new_G4576, new_G7565, new_G7566, new_G7573, new_G7574, new_G4936,
    new_G4937, new_G4977, new_G4978, new_G5105, new_G5359, new_G5362,
    new_G5529, new_G5675, new_G5932, new_G5977, new_G6052, new_G6063,
    new_G6115, new_G6173, new_G6679, new_G6751, new_G6752, new_G6761,
    new_G6762, new_G6795, new_G6796, new_G6805, new_G6806, new_G6931,
    new_G6983, new_G7047, new_G7129, new_G7279, new_G7280, new_G7289,
    new_G7290, new_G7337, new_G7340, new_G7353, new_G7356, new_G7537,
    new_G7538, new_G7547, new_G7548, new_G7581, new_G7582, new_G7591,
    new_G7592, new_G7595, new_G7598, new_G2342, new_G2353, new_G2371,
    new_G2399, new_G2408, new_G2419, new_G2435, new_G2453, new_G2588,
    new_G2599, new_G2617, new_G2642, new_G2654, new_G2675, new_G2700,
    new_G2733, new_G3050, new_G3060, new_G3069, new_G3080, new_G3091,
    new_G3092, new_G3100, new_G3101, new_G3108, new_G3109, new_G3117,
    new_G3120, new_G3121, new_G3282, new_G3294, new_G3313, new_G3343,
    new_G3352, new_G3364, new_G3380, new_G3398, new_G3416, new_G3525,
    new_G3534, new_G3535, new_G3543, new_G3544, new_G3548, new_G3557,
    new_G3558, new_G3566, new_G3567, new_G3844, new_G3855, new_G3873,
    new_G3898, new_G3910, new_G3931, new_G3956, new_G3988, new_G3996,
    new_G4178, new_G4187, new_G4188, new_G4197, new_G4219, new_G4289,
    new_G4290, new_G4298, new_G4299, new_G4306, new_G4307, new_G4315,
    new_G4316, new_G4325, new_G4334, new_G4342, new_G4350, new_G4351,
    new_G4354, new_G4561, new_G4562, new_G4570, new_G4571, new_G4575,
    new_G4584, new_G4585, new_G4593, new_G4594, new_G4938, new_G4979,
    new_G6753, new_G6754, new_G6763, new_G6764, new_G6797, new_G6798,
    new_G6807, new_G6808, new_G7281, new_G7282, new_G7291, new_G7292,
    new_G7539, new_G7540, new_G7549, new_G7550, new_G7583, new_G7584,
    new_G7593, new_G7594, new_G1856, new_G920, new_G925, new_G926,
    new_G927, new_G928, new_G937, new_G938, new_G939, new_G940, new_G941,
    new_G942, new_G943, new_G944, new_G945, new_G946, new_G947, new_G948,
    new_G949, new_G956, new_G1122, new_G1125, new_G1126, new_G1127,
    new_G1128, new_G1132, new_G1133, new_G1134, new_G1137, new_G1138,
    new_G1141, new_G1221, new_G1230, new_G1244, new_G1253, new_G1267,
    new_G1276, new_G1284, new_G1288, new_G1292, new_G1296, new_G1300,
    new_G1304, new_G1702, new_G1705, new_G1706, new_G1707, new_G1709,
    new_G1710, new_G1711, new_G1712, new_G1713, new_G1714, new_G1718,
    new_G1722, new_G1723, new_G1724, new_G1725, new_G1733, new_G1734,
    new_G1735, new_G1736, new_G1737, new_G1738, new_G1739, new_G1740,
    new_G1741, new_G1742, new_G1743, new_G1744, new_G1745, new_G1749,
    new_G1750, new_G1935, new_G1938, new_G1939, new_G1940, new_G1942,
    new_G1943, new_G1944, new_G1945, new_G1946, new_G1947, new_G1948,
    new_G1949, new_G1950, new_G1953, new_G1954, new_G1955, new_G1956,
    new_G1960, new_G1961, new_G1962, new_G1965, new_G1966, new_G1969,
    new_G2343, new_G2354, new_G2372, new_G2400, new_G2409, new_G2420,
    new_G2436, new_G2454, new_G2470, new_G5936, new_G5983, new_G2589,
    new_G2600, new_G2618, new_G2643, new_G2655, new_G2676, new_G2701,
    new_G2734, new_G2740, new_G6056, new_G3022, new_G3025, new_G3026,
    new_G3027, new_G3029, new_G3030, new_G3031, new_G3032, new_G3033,
    new_G3052, new_G3062, new_G3071, new_G3082, new_G3093, new_G3102,
    new_G3110, new_G3119, new_G3122, new_G3228, new_G3231, new_G3232,
    new_G3233, new_G3234, new_G3283, new_G3295, new_G3314, new_G3344,
    new_G3353, new_G3365, new_G3381, new_G3399, new_G3417, new_G6685,
    new_G3508, new_G3517, new_G3527, new_G3536, new_G3545, new_G3550,
    new_G3559, new_G3568, new_G3571, new_G3575, new_G3845, new_G3856,
    new_G3874, new_G3899, new_G3911, new_G3932, new_G3957, new_G3989,
    new_G3997, new_G4180, new_G4189, new_G4198, new_G4207, new_G4216,
    new_G4221, new_G4230, new_G4239, new_G4263, new_G4267, new_G4291,
    new_G4300, new_G4308, new_G4317, new_G4327, new_G4336, new_G4344,
    new_G4352, new_G4355, new_G4535, new_G4544, new_G4558, new_G4563,
    new_G4572, new_G4577, new_G4586, new_G4595, new_G4598, new_G4602,
    new_G4716, new_G4724, new_G4732, new_G4740, new_G4748, new_G4756,
    new_G4764, new_G4772, new_G4780, new_G4788, new_G4939, new_G4980,
    new_G5044, new_G5054, new_G5064, new_G5074, new_G5084, new_G5094,
    new_G5132, new_G5142, new_G5152, new_G5162, new_G5365, new_G5366,
    new_G5488, new_G5498, new_G5508, new_G5518, new_G5546, new_G5556,
    new_G5566, new_G5576, new_G5614, new_G5624, new_G5634, new_G5644,
    new_G5654, new_G5664, new_G5702, new_G5712, new_G5722, new_G5732,
    new_G5820, new_G5828, new_G5836, new_G5844, new_G5852, new_G5860,
    new_G6121, new_G6179, new_G6261, new_G7359, new_G7360, new_G7343,
    new_G7344, new_G6809, new_G6812, new_G6819, new_G6822, new_G6989,
    new_G7135, new_G7345, new_G7348, new_G7601, new_G7602, new_G7603,
    new_G7606, new_G7611, new_G7614, new_G929, new_G950, new_G1129,
    new_G1708, new_G1715, new_G1726, new_G1746, new_G1941, new_G1957,
    new_G2471, new_G2741, new_G3028, new_G3034, new_G3235, new_G5014,
    new_G5034, new_G5102, new_G5122, new_G5367, new_G5368, new_G5478,
    new_G5536, new_G5584, new_G5604, new_G5672, new_G5692, new_G5817,
    new_G5825, new_G5833, new_G5841, new_G6340, new_G6341, new_G6350,
    new_G6351, new_G7436, new_G7437, new_G4720, new_G4728, new_G4736,
    new_G4744, new_G4752, new_G4760, new_G4768, new_G4776, new_G4784,
    new_G4792, new_G3350, new_G2406, new_G924, new_G5088, new_G5098,
    new_G997, new_G1146, new_G1287, new_G1291, new_G1295, new_G1299,
    new_G1303, new_G1307, new_G1309, new_G1312, new_G1315, new_G1318,
    new_G1321, new_G1324, new_G1721, new_G5522, new_G5580, new_G5658,
    new_G5668, new_G1788, new_G1974, new_G5824, new_G5832, new_G5840,
    new_G5848, new_G1999, new_G5856, new_G2003, new_G5864, new_G2472,
    new_G2487, new_G2492, new_G2493, new_G2494, new_G2500, new_G2501,
    new_G2502, new_G2503, new_G2504, new_G2505, new_G2506, new_G2507,
    new_G2511, new_G2512, new_G2513, new_G2514, new_G2518, new_G2519,
    new_G2520, new_G2523, new_G2524, new_G2527, new_G2742, new_G2749,
    new_G2754, new_G2755, new_G2756, new_G2762, new_G2763, new_G2764,
    new_G2765, new_G2766, new_G2767, new_G2776, new_G2777, new_G2778,
    new_G2779, new_G2788, new_G2789, new_G2790, new_G2792, new_G2793,
    new_G2794, new_G2795, new_G2796, new_G2798, new_G2799, new_G2800,
    new_G2804, new_G3035, new_G3045, new_G3123, new_G3128, new_G3129,
    new_G3130, new_G3136, new_G3139, new_G3140, new_G3141, new_G3142,
    new_G3249, new_G3431, new_G3434, new_G3435, new_G3436, new_G3438,
    new_G3439, new_G3440, new_G3441, new_G3442, new_G3443, new_G3444,
    new_G3445, new_G3446, new_G3449, new_G3450, new_G3451, new_G3452,
    new_G3456, new_G3457, new_G3458, new_G3460, new_G3461, new_G3463,
    new_G3531, new_G3540, new_G3554, new_G3563, new_G3574, new_G3578,
    new_G3579, new_G3583, new_G3587, new_G3591, new_G3596, new_G3599,
    new_G4004, new_G4007, new_G4008, new_G4009, new_G4011, new_G4012,
    new_G4013, new_G4014, new_G4015, new_G4016, new_G4020, new_G4024,
    new_G4025, new_G4026, new_G4027, new_G4035, new_G4036, new_G4037,
    new_G4038, new_G4039, new_G4040, new_G4041, new_G4042, new_G4043,
    new_G4044, new_G4045, new_G4046, new_G4047, new_G4051, new_G4052,
    new_G4184, new_G4193, new_G4247, new_G4251, new_G4255, new_G4259,
    new_G4266, new_G4270, new_G4284, new_G4287, new_G4356, new_G4361,
    new_G4362, new_G4363, new_G4369, new_G4372, new_G4373, new_G4374,
    new_G4375, new_G4567, new_G4581, new_G4590, new_G4601, new_G4605,
    new_G4606, new_G4610, new_G4614, new_G4618, new_G4623, new_G4626,
    new_G4796, new_G4804, new_G4812, new_G4820, new_G4828, new_G4844,
    new_G4852, new_G4860, new_G4868, new_G4945, new_G4948, new_G4986,
    new_G4989, new_G5048, new_G5058, new_G5068, new_G5078, new_G5166,
    new_G5136, new_G5146, new_G5156, new_G5388, new_G5492, new_G5502,
    new_G5512, new_G5550, new_G5560, new_G5570, new_G5618, new_G5628,
    new_G5638, new_G5648, new_G5736, new_G5706, new_G5716, new_G5726,
    new_G5940, new_G5948, new_G5956, new_G5964, new_G5972, new_G5980,
    new_G6080, new_G6090, new_G6100, new_G6110, new_G6138, new_G6148,
    new_G6158, new_G6168, new_G6216, new_G6226, new_G6236, new_G6246,
    new_G6256, new_G6267, new_G6304, new_G6314, new_G6324, new_G6342,
    new_G6352, new_G7351, new_G7352, new_G6642, new_G6650, new_G6658,
    new_G6666, new_G6674, new_G6682, new_G6815, new_G6816, new_G6825,
    new_G6826, new_G6948, new_G6958, new_G6968, new_G6978, new_G7006,
    new_G7016, new_G7026, new_G7036, new_G7074, new_G7084, new_G7094,
    new_G7104, new_G7114, new_G7124, new_G7162, new_G7172, new_G7182,
    new_G7192, new_G7438, new_G7617, new_G7618, new_G7609, new_G7610,
    new_G1151, new_G1002, new_G933, new_G1308, new_G1311, new_G1314,
    new_G1317, new_G1320, new_G1323, new_G1730, new_G1789, new_G1981,
    new_G5823, new_G1986, new_G5831, new_G1989, new_G5839, new_G1993,
    new_G5847, new_G1996, new_G2000, new_G2004, new_G2495, new_G2515,
    new_G2757, new_G2768, new_G2780, new_G2801, new_G3046, new_G3131,
    new_G3143, new_G3238, new_G3258, new_G3437, new_G3453, new_G3595,
    new_G3598, new_G4010, new_G4017, new_G4028, new_G4048, new_G4283,
    new_G4286, new_G4364, new_G4376, new_G4622, new_G4625, new_G4947,
    new_G4988, new_G5018, new_G5019, new_G5024, new_G5038, new_G5106,
    new_G5107, new_G5112, new_G5126, new_G5468, new_G5482, new_G5526,
    new_G5540, new_G5588, new_G5589, new_G5594, new_G5608, new_G5676,
    new_G5677, new_G5682, new_G5696, new_G5937, new_G5945, new_G5953,
    new_G5961, new_G6070, new_G6128, new_G6264, new_G6284, new_G6360,
    new_G6361, new_G6639, new_G6647, new_G6655, new_G6663, new_G6817,
    new_G6818, new_G6827, new_G6828, new_G6938, new_G6996, new_G7044,
    new_G7064, new_G7132, new_G7152, new_G7446, new_G7447, new_G7456,
    new_G7457, new_G241, new_G265, new_G2005, new_G4800, new_G4808,
    new_G4816, new_G4824, new_G4832, new_G4848, new_G4856, new_G4864,
    new_G4872, new_G1310, new_G1313, new_G1316, new_G1319, new_G1322,
    new_G1325, new_G5392, new_G1790, new_G1982, new_G1985, new_G1988,
    new_G1992, new_G1995, new_G2001, new_G2491, new_G2508, new_G2522,
    new_G2526, new_G2529, new_G2531, new_G5944, new_G5952, new_G5960,
    new_G5968, new_G2555, new_G5976, new_G2559, new_G5984, new_G2753,
    new_G2771, new_G2791, new_G2797, new_G2807, new_G6114, new_G6172,
    new_G6250, new_G6260, new_G6346, new_G6356, new_G3127, new_G3156,
    new_G3259, new_G3466, new_G6646, new_G6654, new_G6662, new_G6670,
    new_G3483, new_G6678, new_G3487, new_G6686, new_G3582, new_G3586,
    new_G3590, new_G3594, new_G3597, new_G3600, new_G3602, new_G3605,
    new_G3608, new_G3611, new_G4023, new_G6982, new_G7040, new_G7118,
    new_G7128, new_G4089, new_G4250, new_G4254, new_G4258, new_G4262,
    new_G4272, new_G4275, new_G4278, new_G4281, new_G4285, new_G4288,
    new_G4360, new_G4380, new_G4386, new_G7442, new_G4609, new_G4613,
    new_G4617, new_G4621, new_G4624, new_G4627, new_G4629, new_G4632,
    new_G4635, new_G4638, new_G4836, new_G4949, new_G4990, new_G5020,
    new_G5108, new_G5590, new_G5678, new_G6084, new_G6094, new_G6104,
    new_G6142, new_G6152, new_G6162, new_G6206, new_G6220, new_G6230,
    new_G6240, new_G6328, new_G6294, new_G6308, new_G6318, new_G6362,
    new_G6840, new_G6848, new_G6952, new_G6962, new_G6972, new_G7010,
    new_G7020, new_G7030, new_G7078, new_G7088, new_G7098, new_G7108,
    new_G7196, new_G7166, new_G7176, new_G7186, new_G7448, new_G7458,
    new_G254, new_G260, new_G1987, new_G1994, new_G2002, new_G962,
    new_G1751, new_G1990, new_G1997, new_G2499, new_G2536, new_G5943,
    new_G2542, new_G5951, new_G2545, new_G5959, new_G2549, new_G5967,
    new_G2552, new_G2556, new_G2560, new_G2761, new_G2784, new_G2853,
    new_G3135, new_G3146, new_G3163, new_G3467, new_G6645, new_G3470,
    new_G6653, new_G3473, new_G6661, new_G3477, new_G6669, new_G3480,
    new_G3484, new_G3488, new_G3601, new_G3604, new_G3607, new_G3610,
    new_G4032, new_G4090, new_G4271, new_G4274, new_G4277, new_G4280,
    new_G4368, new_G4379, new_G4387, new_G4628, new_G4631, new_G4634,
    new_G4637, new_G4841, new_G4849, new_G4857, new_G4865, new_G5021,
    new_G5028, new_G5109, new_G5116, new_G5369, new_G5377, new_G5385,
    new_G5472, new_G5473, new_G5530, new_G5531, new_G5591, new_G5598,
    new_G5679, new_G5686, new_G6060, new_G6074, new_G6118, new_G6132,
    new_G6176, new_G6186, new_G6196, new_G6268, new_G6269, new_G6274,
    new_G6288, new_G6337, new_G6829, new_G6928, new_G6942, new_G6986,
    new_G7000, new_G7048, new_G7049, new_G7054, new_G7068, new_G7136,
    new_G7137, new_G7142, new_G7156, new_G7433, new_G242, new_G3151,
    new_G257, new_G263, new_G266, new_G1991, new_G1998, new_G3489,
    new_G371, new_G4840, new_G2561, new_G2532, new_G2537, new_G2541,
    new_G2544, new_G2548, new_G2551, new_G2557, new_G2563, new_G2577,
    new_G2775, new_G2806, new_G2808, new_G2852, new_G2854, new_G6366,
    new_G4381, new_G3164, new_G3241, new_G3468, new_G3469, new_G3472,
    new_G3476, new_G3479, new_G3485, new_G3603, new_G3606, new_G3609,
    new_G3612, new_G6844, new_G6852, new_G4091, new_G4273, new_G4276,
    new_G4279, new_G4282, new_G4382, new_G4388, new_G7452, new_G7462,
    new_G4630, new_G4633, new_G4636, new_G4639, new_G4955, new_G4958,
    new_G4996, new_G4999, new_G5474, new_G5532, new_G6210, new_G6270,
    new_G6298, new_G7050, new_G7138, new_G3471, new_G3478, new_G3486,
    new_G372, new_G2543, new_G2550, new_G2558, new_G4847, new_G387,
    new_G4855, new_G390, new_G4863, new_G393, new_G4871, new_G396,
    new_G965, new_G5375, new_G1327, new_G5383, new_G1330, new_G5391,
    new_G1333, new_G1754, new_G2546, new_G2553, new_G2564, new_G2809,
    new_G2813, new_G6345, new_G2860, new_G3474, new_G3481, new_G6835,
    new_G3614, new_G4053, new_G7441, new_G4516, new_G4957, new_G4998,
    new_G5027, new_G5030, new_G5115, new_G5118, new_G5475, new_G5533,
    new_G5597, new_G5600, new_G5685, new_G5688, new_G6064, new_G6065,
    new_G6122, new_G6123, new_G6180, new_G6181, new_G6190, new_G6200,
    new_G6271, new_G6278, new_G6347, new_G6357, new_G6837, new_G6845,
    new_G6932, new_G6933, new_G6990, new_G6991, new_G7051, new_G7058,
    new_G7139, new_G7146, new_G7443, new_G7453, new_G243, new_G244,
    new_G245, new_G255, new_G256, new_G261, new_G262, new_G267, new_G268,
    new_G269, new_G3475, new_G3482, new_G2547, new_G2554, new_G386,
    new_G389, new_G392, new_G395, new_G1326, new_G1329, new_G1332,
    new_G1436, new_G1440, new_G1445, new_G1450, new_G1454, new_G2859,
    new_G4385, new_G3148, new_G3239, new_G3240, new_G3265, new_G3267,
    new_G3270, new_G3274, new_G3277, new_G3613, new_G4515, new_G4959,
    new_G5000, new_G5029, new_G5117, new_G5599, new_G5687, new_G6066,
    new_G6124, new_G6182, new_G6934, new_G6992, new_G375, new_G378,
    new_G381, new_G384, new_G1328, new_G1331, new_G1334, new_G1447,
    new_G1766, new_G2571, new_G2579, new_G2812, new_G2816, new_G2851,
    new_G2861, new_G6355, new_G2863, new_G6365, new_G2866, new_G3147,
    new_G3242, new_G3271, new_G3279, new_G3615, new_G6843, new_G3617,
    new_G6851, new_G3620, new_G4056, new_G4517, new_G7451, new_G4519,
    new_G7461, new_G4522, new_G5031, new_G5119, new_G5481, new_G5484,
    new_G5539, new_G5542, new_G5601, new_G5689, new_G6067, new_G6125,
    new_G6183, new_G6277, new_G6280, new_G6935, new_G6993, new_G7057,
    new_G7060, new_G7145, new_G7148, new_G4968, new_G5009, new_G2850,
    new_G2862, new_G2865, new_G3149, new_G3243, new_G3616, new_G3619,
    new_G4518, new_G4521, new_G4965, new_G5006, new_G5483, new_G5541,
    new_G6279, new_G7059, new_G7147, new_G374, new_G377, new_G380,
    new_G383, new_G955, new_G4967, new_G5008, new_G975, new_G1136,
    new_G1140, new_G1143, new_G1145, new_G1160, new_G1771, new_G1964,
    new_G1968, new_G1971, new_G1973, new_G2007, new_G2578, new_G2864,
    new_G2867, new_G3150, new_G3245, new_G3618, new_G3621, new_G4067,
    new_G4520, new_G4523, new_G4713, new_G4753, new_G5037, new_G5040,
    new_G5125, new_G5128, new_G5485, new_G5543, new_G5607, new_G5610,
    new_G5695, new_G5698, new_G6073, new_G6076, new_G6131, new_G6134,
    new_G6189, new_G6192, new_G6281, new_G6941, new_G6944, new_G6999,
    new_G7002, new_G7061, new_G7149, new_G958, new_G967, new_G971,
    new_G1161, new_G2008, new_G2580, new_G2868, new_G3152, new_G4443,
    new_G4524, new_G4721, new_G4729, new_G4737, new_G4745, new_G4761,
    new_G4769, new_G4777, new_G4785, new_G5039, new_G5127, new_G5609,
    new_G5697, new_G6075, new_G6133, new_G6191, new_G6943, new_G7001,
    new_G3248, new_G248, new_G4719, new_G294, new_G4759, new_G323,
    new_G980, new_G4072, new_G5041, new_G5129, new_G5491, new_G5494,
    new_G5549, new_G5552, new_G5611, new_G5699, new_G6077, new_G6135,
    new_G6193, new_G6287, new_G6290, new_G6945, new_G7003, new_G7067,
    new_G7070, new_G7155, new_G7158, new_G247, new_G3155, new_G251,
    new_G272, new_G961, new_G275, new_G293, new_G297, new_G300, new_G303,
    new_G306, new_G4727, new_G309, new_G4735, new_G312, new_G4743,
    new_G315, new_G4751, new_G318, new_G322, new_G4767, new_G326,
    new_G4775, new_G329, new_G4783, new_G332, new_G4791, new_G335,
    new_G2881, new_G993, new_G994, new_G1166, new_G1171, new_G1174,
    new_G2014, new_G3459, new_G3462, new_G3464, new_G3465, new_G3490,
    new_G4793, new_G5493, new_G5551, new_G6289, new_G7069, new_G7157,
    new_G250, new_G274, new_G308, new_G311, new_G314, new_G317, new_G325,
    new_G328, new_G331, new_G334, new_G417, new_G991, new_G992, new_G3491,
    new_G4801, new_G4809, new_G4817, new_G4825, new_G5047, new_G5050,
    new_G5135, new_G5138, new_G5495, new_G5553, new_G5617, new_G5620,
    new_G5705, new_G5708, new_G6083, new_G6086, new_G6141, new_G6144,
    new_G6199, new_G6202, new_G6291, new_G6951, new_G6954, new_G7009,
    new_G7012, new_G7071, new_G7159, new_G271, new_G296, new_G299,
    new_G302, new_G305, new_G4799, new_G343, new_G1170, new_G1173,
    new_G5049, new_G5137, new_G5167, new_G5619, new_G5707, new_G6085,
    new_G6143, new_G6201, new_G6953, new_G7011, new_G342, new_G346,
    new_G349, new_G352, new_G355, new_G4807, new_G358, new_G4815, new_G361,
    new_G4823, new_G364, new_G4831, new_G367, new_G1172, new_G1175,
    new_G3497, new_G5051, new_G5139, new_G5501, new_G5504, new_G5559,
    new_G5562, new_G5621, new_G5709, new_G6087, new_G6145, new_G6203,
    new_G6297, new_G6300, new_G6955, new_G7013, new_G7077, new_G7080,
    new_G7165, new_G7168, new_G357, new_G360, new_G363, new_G366,
    new_G5173, new_G5503, new_G5561, new_G6299, new_G7079, new_G7167,
    new_G345, new_G348, new_G351, new_G354, new_G5057, new_G5060,
    new_G5145, new_G5148, new_G5505, new_G5563, new_G5627, new_G5630,
    new_G5715, new_G5718, new_G6093, new_G6096, new_G6151, new_G6154,
    new_G6209, new_G6212, new_G6301, new_G6961, new_G6964, new_G7019,
    new_G7022, new_G7081, new_G7169, new_G5059, new_G5147, new_G5629,
    new_G5717, new_G6095, new_G6153, new_G6211, new_G6963, new_G7021,
    new_G5061, new_G5149, new_G5511, new_G5514, new_G5569, new_G5572,
    new_G5631, new_G5719, new_G6097, new_G6155, new_G6213, new_G6307,
    new_G6310, new_G6965, new_G7023, new_G7087, new_G7090, new_G7175,
    new_G7178, new_G5513, new_G5571, new_G6309, new_G7089, new_G7177,
    new_G5067, new_G5070, new_G5155, new_G5158, new_G5515, new_G5573,
    new_G5637, new_G5640, new_G5725, new_G5728, new_G6103, new_G6106,
    new_G6161, new_G6164, new_G6219, new_G6222, new_G6311, new_G6971,
    new_G6974, new_G7029, new_G7032, new_G7091, new_G7179, new_G5069,
    new_G5157, new_G5639, new_G5727, new_G6105, new_G6163, new_G6221,
    new_G6973, new_G7031, new_G5521, new_G1756, new_G5579, new_G1761,
    new_G5071, new_G5159, new_G5641, new_G5729, new_G6107, new_G6165,
    new_G6223, new_G6317, new_G6320, new_G6975, new_G7033, new_G7097,
    new_G7100, new_G7185, new_G7188, new_G1755, new_G1760, new_G6319,
    new_G7099, new_G7187, new_G1757, new_G1762, new_G6113, new_G2818,
    new_G6171, new_G2823, new_G6981, new_G4058, new_G7039, new_G4063,
    new_G5077, new_G5080, new_G5165, new_G5090, new_G5647, new_G5650,
    new_G5735, new_G5660, new_G6229, new_G6232, new_G6321, new_G7101,
    new_G7189, new_G2817, new_G2822, new_G4057, new_G4062, new_G5079,
    new_G5089, new_G5649, new_G5659, new_G6231, new_G1782, new_G1783,
    new_G1784, new_G1785, new_G2819, new_G2824, new_G4059, new_G4064,
    new_G5081, new_G5091, new_G5651, new_G5661, new_G6233, new_G6327,
    new_G6252, new_G7107, new_G7110, new_G7195, new_G7120, new_G5737,
    new_G6251, new_G7109, new_G7119, new_G5087, new_G985, new_G5097,
    new_G988, new_G5657, new_G1776, new_G5667, new_G1779, new_G2844,
    new_G2845, new_G2846, new_G2847, new_G4083, new_G4084, new_G4085,
    new_G4086, new_G6239, new_G6242, new_G6253, new_G7111, new_G7121,
    new_G984, new_G987, new_G1775, new_G1778, new_G5743, new_G6241,
    new_G6329, new_G7197, new_G986, new_G989, new_G1777, new_G1780,
    new_G6259, new_G2841, new_G7117, new_G4077, new_G7127, new_G4080,
    new_G6243, new_G990, new_G996, new_G1781, new_G1787, new_G2840,
    new_G6335, new_G4076, new_G4079, new_G7203, new_G995, new_G1786,
    new_G6249, new_G2838, new_G2842, new_G4078, new_G4081, new_G2837,
    new_G2843, new_G4082, new_G4088, new_G5170, new_G5740, new_G2839,
    new_G2848, new_G4087, new_G1791, new_G1003, new_G5174, new_G5744,
    new_G2849, new_G7200, new_G1792, new_G1004, new_G6332, new_G320,
    new_G337, new_G4092, new_G7204, new_G4093, new_G2855, new_G6336,
    new_G369, new_G2856, new_G398;
  assign G2 = G1;
  assign G3 = G1;
  assign new_G400 = ~G57;
  assign new_G1184 = G134 & G133;
  assign G450 = G1459;
  assign G448 = G1469;
  assign G444 = G1480;
  assign G442 = G1486;
  assign G440 = G1492;
  assign G438 = G1496;
  assign new_G1501 = G199 & G188 & G162 & G172;
  assign G496 = G2208;
  assign G494 = G2218;
  assign G492 = G2224;
  assign G490 = G2230;
  assign G488 = G2236;
  assign G486 = G2239;
  assign G484 = G2247;
  assign G482 = G2253;
  assign G480 = G2256;
  assign new_G2857 = G240 & G228 & G150 & G184;
  assign G560 = G3698;
  assign G542 = G3701;
  assign G558 = G3705;
  assign G556 = G3711;
  assign G554 = G3717;
  assign G552 = G3723;
  assign G550 = G3729;
  assign G548 = G3737;
  assign G546 = G3743;
  assign G544 = G3749;
  assign G540 = G4393;
  assign G538 = G4400;
  assign G536 = G4405;
  assign G534 = G4410;
  assign G532 = G4415;
  assign G530 = G4420;
  assign G528 = G4427;
  assign G526 = G4432;
  assign G524 = G4437;
  assign new_G4442 = G186 & G185 & G183 & G182;
  assign new_G4514 = G230 & G218 & G210 & G152;
  assign G279 = ~G15;
  assign new_G401 = ~G5;
  assign new_G573 = G1;
  assign new_G574 = ~G5;
  assign new_G575 = ~G5;
  assign new_G1178 = ~G2236;
  assign new_G1186 = ~G2253;
  assign new_G1192 = ~G2256;
  assign new_G1198 = G38;
  assign new_G1205 = G15;
  assign new_G1206 = ~G12 | ~G9;
  assign new_G1207 = ~G12 | ~G9;
  assign new_G1210 = G38;
  assign new_G1458 = ~G1455;
  assign new_G1461 = ~G1459;
  assign G436 = G1462;
  assign new_G1464 = ~G1462;
  assign new_G1471 = ~G1469;
  assign new_G1475 = G106;
  assign new_G1482 = ~G1480;
  assign new_G1488 = ~G1486;
  assign new_G1495 = ~G1492;
  assign new_G1499 = ~G1496;
  assign new_G1500 = ~G106;
  assign new_G1503 = G18;
  assign new_G1512 = G18;
  assign new_G1518 = G4528 & G1492;
  assign new_G1524 = G18;
  assign new_G1535 = ~G18;
  assign new_G1541 = ~G4528 | ~G1496;
  assign new_G2207 = ~G2204;
  assign new_G2210 = ~G2208;
  assign G478 = G2211;
  assign new_G2213 = ~G2211;
  assign new_G2220 = ~G2218;
  assign new_G2226 = ~G2224;
  assign new_G2232 = ~G2230;
  assign new_G2238 = ~G2236;
  assign new_G2241 = ~G2239;
  assign new_G2249 = ~G2247;
  assign new_G2255 = ~G2253;
  assign new_G2258 = ~G2256;
  assign new_G2828 = G4526;
  assign new_G3700 = ~G3698;
  assign new_G3703 = ~G3701;
  assign new_G3707 = ~G3705;
  assign new_G3713 = ~G3711;
  assign new_G3719 = ~G3717;
  assign new_G3725 = ~G3723;
  assign new_G3731 = ~G3729;
  assign new_G3739 = ~G3737;
  assign new_G3745 = ~G3743;
  assign new_G3751 = ~G3749;
  assign new_G4121 = ~G4393;
  assign G522 = G4394;
  assign new_G4396 = ~G4394;
  assign new_G4402 = ~G4400;
  assign new_G4407 = ~G4405;
  assign new_G4412 = ~G4410;
  assign new_G4417 = ~G4415;
  assign new_G4422 = ~G4420;
  assign new_G4429 = ~G4427;
  assign new_G4434 = ~G4432;
  assign new_G4439 = ~G4437;
  assign new_G4833 = G4526;
  assign G402 = ~new_G400 | ~new_G401;
  assign G404 = ~new_G2857;
  assign G406 = ~new_G4514;
  assign G408 = ~new_G4442;
  assign G410 = ~new_G1501;
  assign new_G2876 = new_G2857 & new_G4514;
  assign new_G2878 = new_G4442 & new_G1501;
  assign G432 = new_G573;
  assign G446 = new_G1475;
  assign new_G1519 = ~new_G1518;
  assign new_G2871 = G4528 & new_G1458;
  assign new_G2883 = ~G4528 | ~new_G2207;
  assign new_G280 = new_G1184 & new_G575;
  assign G284 = ~G1197 | ~new_G574;
  assign G286 = ~new_G1205;
  assign G289 = ~G1197 | ~new_G574;
  assign G292 = ~new_G1184 | ~new_G575;
  assign G341 = ~new_G1205;
  assign new_G4839 = ~new_G4833;
  assign new_G572 = new_G573;
  assign new_G581 = new_G1206;
  assign new_G587 = new_G1512;
  assign new_G601 = new_G1206;
  assign new_G606 = new_G1512;
  assign new_G650 = new_G1206;
  assign new_G657 = new_G1512;
  assign new_G671 = new_G1207;
  assign new_G678 = new_G1503;
  assign new_G777 = new_G1541 & new_G1198;
  assign new_G1115 = new_G1541 & new_G1198;
  assign new_G1336 = new_G1512;
  assign new_G1350 = new_G1503;
  assign new_G1477 = ~new_G1475;
  assign new_G1507 = ~new_G1503;
  assign new_G1514 = ~new_G1512;
  assign new_G1530 = ~new_G1524;
  assign new_G2259 = new_G1535;
  assign new_G2833 = ~new_G2828;
  assign new_G2872 = ~new_G2871;
  assign new_G2886 = new_G1207;
  assign new_G2892 = new_G1503;
  assign new_G2905 = new_G1207;
  assign new_G2909 = new_G1503;
  assign new_G3622 = new_G1524;
  assign new_G3635 = new_G1524;
  assign new_G3755 = new_G1535;
  assign new_G4640 = new_G1524;
  assign new_G4653 = new_G1524;
  assign new_G4873 = new_G1541;
  assign new_G4876 = new_G1198;
  assign new_G4881 = new_G1488;
  assign new_G4889 = new_G1482;
  assign new_G4905 = new_G1471;
  assign new_G4916 = new_G1198;
  assign new_G4921 = new_G1464;
  assign new_G5175 = new_G1541;
  assign new_G5178 = new_G1198;
  assign new_G5186 = new_G1198;
  assign new_G5191 = new_G1488;
  assign new_G5199 = new_G1482;
  assign new_G5215 = new_G1471;
  assign new_G5223 = new_G1464;
  assign new_G5393 = new_G1192;
  assign new_G5401 = new_G1186;
  assign new_G5409 = new_G2249;
  assign new_G5417 = new_G1178;
  assign new_G5425 = new_G2232;
  assign new_G5433 = new_G2226;
  assign new_G5441 = new_G2220;
  assign new_G5449 = new_G2241;
  assign new_G5457 = new_G2213;
  assign new_G5745 = new_G1192;
  assign new_G5753 = new_G1186;
  assign new_G5761 = new_G2249;
  assign new_G5769 = new_G2241;
  assign new_G5777 = new_G1178;
  assign new_G5785 = new_G2232;
  assign new_G5793 = new_G2226;
  assign new_G5801 = new_G2220;
  assign new_G5809 = new_G2213;
  assign new_G5865 = new_G3751;
  assign new_G5873 = new_G3745;
  assign new_G5881 = new_G3739;
  assign new_G5889 = new_G3731;
  assign new_G5897 = new_G3725;
  assign new_G5905 = new_G3719;
  assign new_G5913 = new_G3713;
  assign new_G5921 = new_G3707;
  assign new_G5985 = new_G3751;
  assign new_G5993 = new_G3745;
  assign new_G6001 = new_G3739;
  assign new_G6009 = new_G3725;
  assign new_G6017 = new_G3719;
  assign new_G6025 = new_G3713;
  assign new_G6033 = new_G3707;
  assign new_G6041 = new_G3731;
  assign new_G6514 = new_G1210;
  assign new_G6554 = new_G1210;
  assign new_G6567 = new_G4439;
  assign new_G6575 = new_G4434;
  assign new_G6583 = new_G4429;
  assign new_G6591 = new_G4422;
  assign new_G6599 = new_G4417;
  assign new_G6607 = new_G4412;
  assign new_G6615 = new_G4407;
  assign new_G6623 = new_G4402;
  assign new_G6631 = new_G4396;
  assign new_G6853 = new_G4439;
  assign new_G6861 = new_G4434;
  assign new_G6869 = new_G4429;
  assign new_G6877 = new_G4417;
  assign new_G6885 = new_G4412;
  assign new_G6893 = new_G4407;
  assign new_G6901 = new_G4402;
  assign new_G6909 = new_G4422;
  assign new_G6917 = new_G4396;
  assign G281 = ~new_G280;
  assign G453 = new_G572;
  assign new_G784 = new_G1519 & new_G1198;
  assign new_G1014 = new_G1198 & new_G1519;
  assign new_G3221 = new_G2883 & new_G1210;
  assign new_G4913 = new_G1519;
  assign new_G4929 = ~new_G1519 & ~new_G1198;
  assign new_G5183 = new_G1519;
  assign new_G5231 = ~new_G1198 & ~new_G1519;
  assign new_G6511 = new_G2883;
  assign G278 = G163 & new_G572;
  assign new_G615 = G170 & new_G587;
  assign new_G594 = ~new_G587;
  assign new_G611 = ~new_G606;
  assign new_G617 = G169 & new_G587;
  assign new_G619 = G168 & new_G587;
  assign new_G621 = G167 & new_G587;
  assign new_G623 = G166 & new_G606;
  assign new_G625 = G165 & new_G606;
  assign new_G627 = G164 & new_G606;
  assign new_G664 = ~new_G657;
  assign new_G685 = ~new_G678;
  assign new_G691 = G177 & new_G657;
  assign new_G693 = G176 & new_G657;
  assign new_G695 = G175 & new_G657;
  assign new_G697 = G174 & new_G657;
  assign new_G699 = G173 & new_G657;
  assign new_G701 = G157 & new_G678;
  assign new_G703 = G156 & new_G678;
  assign new_G705 = G155 & new_G678;
  assign new_G707 = G154 & new_G678;
  assign new_G709 = G153 & new_G678;
  assign new_G4879 = ~new_G4873;
  assign new_G4880 = ~new_G4876;
  assign new_G4887 = ~new_G4881;
  assign new_G4895 = ~new_G4889;
  assign new_G4911 = ~new_G4905;
  assign new_G4920 = ~new_G4916;
  assign new_G4927 = ~new_G4921;
  assign new_G5181 = ~new_G5175;
  assign new_G5182 = ~new_G5178;
  assign new_G5190 = ~new_G5186;
  assign new_G5197 = ~new_G5191;
  assign new_G5205 = ~new_G5199;
  assign new_G5221 = ~new_G5215;
  assign new_G5229 = ~new_G5223;
  assign new_G1343 = ~new_G1336;
  assign new_G1357 = ~new_G1350;
  assign new_G1364 = G181 & new_G1336;
  assign new_G1366 = G171 & new_G1336;
  assign new_G1368 = G180 & new_G1336;
  assign new_G1370 = G179 & new_G1336;
  assign new_G1372 = G178 & new_G1336;
  assign new_G1374 = G161 & new_G1350;
  assign new_G1376 = G151 & new_G1350;
  assign new_G1378 = G160 & new_G1350;
  assign new_G1380 = G159 & new_G1350;
  assign new_G1382 = G158 & new_G1350;
  assign new_G5399 = ~new_G5393;
  assign new_G5407 = ~new_G5401;
  assign new_G5415 = ~new_G5409;
  assign new_G5423 = ~new_G5417;
  assign new_G5431 = ~new_G5425;
  assign new_G5439 = ~new_G5433;
  assign new_G5447 = ~new_G5441;
  assign new_G5455 = ~new_G5449;
  assign new_G5463 = ~new_G5457;
  assign new_G5751 = ~new_G5745;
  assign new_G5759 = ~new_G5753;
  assign new_G5767 = ~new_G5761;
  assign new_G5775 = ~new_G5769;
  assign new_G5783 = ~new_G5777;
  assign new_G5791 = ~new_G5785;
  assign new_G5799 = ~new_G5793;
  assign new_G5807 = ~new_G5801;
  assign new_G5815 = ~new_G5809;
  assign new_G2019 = new_G1514;
  assign new_G2032 = new_G1507;
  assign new_G2117 = new_G1514;
  assign new_G2130 = new_G1507;
  assign new_G2266 = ~new_G2259;
  assign new_G2272 = new_G1507;
  assign new_G2286 = G44 & new_G2259;
  assign new_G2288 = G41 & new_G2259;
  assign new_G2290 = G29 & new_G2259;
  assign new_G2292 = G26 & new_G2259;
  assign new_G2294 = G23 & new_G2259;
  assign new_G5871 = ~new_G5865;
  assign new_G5879 = ~new_G5873;
  assign new_G5887 = ~new_G5881;
  assign new_G5895 = ~new_G5889;
  assign new_G5903 = ~new_G5897;
  assign new_G5911 = ~new_G5905;
  assign new_G5919 = ~new_G5913;
  assign new_G5927 = ~new_G5921;
  assign new_G5991 = ~new_G5985;
  assign new_G5999 = ~new_G5993;
  assign new_G6007 = ~new_G6001;
  assign new_G6015 = ~new_G6009;
  assign new_G6023 = ~new_G6017;
  assign new_G6031 = ~new_G6025;
  assign new_G6039 = ~new_G6033;
  assign new_G6047 = ~new_G6041;
  assign new_G2899 = ~new_G2892;
  assign new_G2914 = ~new_G2909;
  assign new_G2919 = G209 & new_G2892;
  assign new_G2921 = G216 & new_G2892;
  assign new_G2923 = G215 & new_G2892;
  assign new_G2925 = G214 & new_G2892;
  assign new_G2927 = G213 & new_G2909;
  assign new_G2929 = G212 & new_G2909;
  assign new_G2931 = G211 & new_G2909;
  assign new_G6518 = ~new_G6514;
  assign new_G3173 = new_G2872 & new_G1210;
  assign new_G6558 = ~new_G6554;
  assign new_G6573 = ~new_G6567;
  assign new_G6581 = ~new_G6575;
  assign new_G6589 = ~new_G6583;
  assign new_G6597 = ~new_G6591;
  assign new_G6605 = ~new_G6599;
  assign new_G6613 = ~new_G6607;
  assign new_G6621 = ~new_G6615;
  assign new_G6629 = ~new_G6623;
  assign new_G6637 = ~new_G6631;
  assign new_G3629 = ~new_G3622;
  assign new_G3642 = ~new_G3635;
  assign new_G3649 = new_G1461 & new_G3622;
  assign new_G3651 = new_G1464 & new_G3622;
  assign new_G3653 = new_G1471 & new_G3622;
  assign new_G3655 = new_G1500 & new_G3622;
  assign new_G3657 = new_G1482 & new_G3622;
  assign new_G3659 = new_G1488 & new_G3635;
  assign new_G3661 = new_G1495 & new_G3635;
  assign new_G3663 = new_G1499 & new_G3635;
  assign new_G3762 = ~new_G3755;
  assign new_G3768 = new_G1507;
  assign new_G3782 = G47 & new_G3755;
  assign new_G3784 = G35 & new_G3755;
  assign new_G3786 = G32 & new_G3755;
  assign new_G3788 = G50 & new_G3755;
  assign new_G3790 = G66 & new_G3755;
  assign new_G6859 = ~new_G6853;
  assign new_G6867 = ~new_G6861;
  assign new_G6875 = ~new_G6869;
  assign new_G6883 = ~new_G6877;
  assign new_G6891 = ~new_G6885;
  assign new_G6899 = ~new_G6893;
  assign new_G6907 = ~new_G6901;
  assign new_G6915 = ~new_G6909;
  assign new_G6923 = ~new_G6917;
  assign new_G4094 = new_G1530;
  assign new_G4107 = new_G1530;
  assign new_G4444 = new_G1530;
  assign new_G4457 = new_G1530;
  assign new_G4647 = ~new_G4640;
  assign new_G4660 = ~new_G4653;
  assign new_G4667 = new_G2210 & new_G4640;
  assign new_G4669 = new_G2213 & new_G4640;
  assign new_G4671 = new_G2220 & new_G4640;
  assign new_G4673 = new_G2226 & new_G4640;
  assign new_G4675 = new_G2232 & new_G4640;
  assign new_G4677 = new_G2238 & new_G4653;
  assign new_G4679 = new_G2241 & new_G4653;
  assign new_G4681 = new_G2249 & new_G4653;
  assign new_G4683 = new_G2255 & new_G4653;
  assign new_G4685 = new_G2258 & new_G4653;
  assign new_G4897 = new_G1477;
  assign new_G5207 = new_G1477;
  assign new_G6551 = new_G2872;
  assign new_G763 = ~new_G4876 | ~new_G4879;
  assign new_G764 = ~new_G4873 | ~new_G4880;
  assign new_G4919 = ~new_G4913;
  assign new_G886 = ~new_G4913 | ~new_G4920;
  assign new_G1005 = ~new_G5178 | ~new_G5181;
  assign new_G1006 = ~new_G5175 | ~new_G5182;
  assign new_G5189 = ~new_G5183;
  assign new_G1018 = ~new_G5183 | ~new_G5190;
  assign new_G5237 = ~new_G5231;
  assign new_G6517 = ~new_G6511;
  assign new_G3169 = ~new_G6511 | ~new_G6518;
  assign new_G4935 = ~new_G4929;
  assign new_G4970 = new_G784;
  assign new_G5239 = new_G1014;
  assign new_G577 = new_G594 | new_G615;
  assign new_G616 = new_G594 | new_G587;
  assign new_G618 = new_G594 | new_G617;
  assign new_G620 = new_G594 | new_G619;
  assign new_G622 = new_G594 | new_G621;
  assign new_G624 = new_G611 | new_G623;
  assign new_G626 = new_G611 | new_G625;
  assign new_G628 = new_G611 | new_G627;
  assign new_G692 = new_G664 | new_G691;
  assign new_G694 = new_G664 | new_G693;
  assign new_G696 = new_G664 | new_G695;
  assign new_G698 = new_G664 | new_G697;
  assign new_G700 = new_G664 | new_G699;
  assign new_G702 = new_G685 | new_G701;
  assign new_G704 = new_G685 | new_G703;
  assign new_G706 = new_G685 | new_G705;
  assign new_G708 = new_G685 | new_G707;
  assign new_G710 = new_G685 | new_G709;
  assign new_G765 = ~new_G763 | ~new_G764;
  assign new_G4903 = ~new_G4897;
  assign new_G885 = ~new_G4916 | ~new_G4919;
  assign new_G1007 = ~new_G1005 | ~new_G1006;
  assign new_G1017 = ~new_G5186 | ~new_G5189;
  assign new_G5213 = ~new_G5207;
  assign new_G1363 = G141 & new_G1343;
  assign new_G1365 = G147 & new_G1343;
  assign new_G1367 = G138 & new_G1343;
  assign new_G1369 = G144 & new_G1343;
  assign new_G1371 = G135 & new_G1343;
  assign new_G1373 = G141 & new_G1357;
  assign new_G1375 = G147 & new_G1357;
  assign new_G1377 = G138 & new_G1357;
  assign new_G1379 = G144 & new_G1357;
  assign new_G1381 = G135 & new_G1357;
  assign new_G2026 = ~new_G2019;
  assign new_G2039 = ~new_G2032;
  assign new_G2046 = G103 & new_G2019;
  assign new_G2048 = G130 & new_G2019;
  assign new_G2050 = G127 & new_G2019;
  assign new_G2052 = G124 & new_G2019;
  assign new_G2054 = G100 & new_G2019;
  assign new_G2056 = G103 & new_G2032;
  assign new_G2058 = G130 & new_G2032;
  assign new_G2060 = G127 & new_G2032;
  assign new_G2062 = G124 & new_G2032;
  assign new_G2064 = G100 & new_G2032;
  assign new_G2124 = ~new_G2117;
  assign new_G2137 = ~new_G2130;
  assign new_G2144 = G115 & new_G2117;
  assign new_G2146 = G118 & new_G2117;
  assign new_G2148 = G97 & new_G2117;
  assign new_G2150 = G94 & new_G2117;
  assign new_G2152 = G121 & new_G2117;
  assign new_G2154 = G115 & new_G2130;
  assign new_G2156 = G118 & new_G2130;
  assign new_G2158 = G97 & new_G2130;
  assign new_G2160 = G94 & new_G2130;
  assign new_G2162 = G121 & new_G2130;
  assign new_G2279 = ~new_G2272;
  assign new_G2285 = G208 & new_G2266;
  assign new_G2287 = G198 & new_G2266;
  assign new_G2289 = G207 & new_G2266;
  assign new_G2291 = G206 & new_G2266;
  assign new_G2293 = G205 & new_G2266;
  assign new_G2296 = G44 & new_G2272;
  assign new_G2298 = G41 & new_G2272;
  assign new_G2300 = G29 & new_G2272;
  assign new_G2302 = G26 & new_G2272;
  assign new_G2304 = G23 & new_G2272;
  assign new_G2918 = new_G2899 | new_G2892;
  assign new_G2920 = new_G2899 | new_G2919;
  assign new_G2922 = new_G2899 | new_G2921;
  assign new_G2924 = new_G2899 | new_G2923;
  assign new_G2926 = new_G2899 | new_G2925;
  assign new_G2928 = new_G2914 | new_G2927;
  assign new_G2930 = new_G2914 | new_G2929;
  assign new_G2932 = new_G2914 | new_G2931;
  assign new_G3168 = ~new_G6514 | ~new_G6517;
  assign new_G6557 = ~new_G6551;
  assign new_G3211 = ~new_G6551 | ~new_G6558;
  assign new_G3648 = G114 & new_G3629;
  assign new_G3650 = G113 & new_G3629;
  assign new_G3652 = G111 & new_G3629;
  assign new_G3654 = G87 & new_G3629;
  assign new_G3656 = G112 & new_G3629;
  assign new_G3658 = G88 & new_G3642;
  assign new_G3660 = G1455 & new_G3642;
  assign new_G3662 = G2204 & new_G3642;
  assign new_G3665 = new_G3703 & new_G3642;
  assign new_G3666 = G70 & new_G3642;
  assign new_G3775 = ~new_G3768;
  assign new_G3781 = G193 & new_G3762;
  assign new_G3783 = G192 & new_G3762;
  assign new_G3785 = G191 & new_G3762;
  assign new_G3787 = G190 & new_G3762;
  assign new_G3789 = G189 & new_G3762;
  assign new_G3792 = G47 & new_G3768;
  assign new_G3794 = G35 & new_G3768;
  assign new_G3796 = G32 & new_G3768;
  assign new_G3798 = G50 & new_G3768;
  assign new_G3800 = G66 & new_G3768;
  assign new_G4101 = ~new_G4094;
  assign new_G4114 = ~new_G4107;
  assign new_G4123 = G58 & new_G4094;
  assign new_G4126 = G77 & new_G4094;
  assign new_G4129 = G78 & new_G4094;
  assign new_G4132 = G59 & new_G4094;
  assign new_G4135 = G81 & new_G4094;
  assign new_G4138 = G80 & new_G4107;
  assign new_G4141 = G79 & new_G4107;
  assign new_G4144 = G60 & new_G4107;
  assign new_G4147 = G61 & new_G4107;
  assign new_G4150 = G62 & new_G4107;
  assign new_G4451 = ~new_G4444;
  assign new_G4464 = ~new_G4457;
  assign new_G4471 = G69 & new_G4444;
  assign new_G4473 = G70 & new_G4444;
  assign new_G4475 = G74 & new_G4444;
  assign new_G4477 = G76 & new_G4444;
  assign new_G4479 = G75 & new_G4444;
  assign new_G4481 = G73 & new_G4457;
  assign new_G4483 = G53 & new_G4457;
  assign new_G4485 = G54 & new_G4457;
  assign new_G4487 = G55 & new_G4457;
  assign new_G4489 = G56 & new_G4457;
  assign new_G4666 = G82 & new_G4647;
  assign new_G4668 = G65 & new_G4647;
  assign new_G4670 = G83 & new_G4647;
  assign new_G4672 = G84 & new_G4647;
  assign new_G4674 = G85 & new_G4647;
  assign new_G4676 = G64 & new_G4660;
  assign new_G4678 = G63 & new_G4660;
  assign new_G4680 = G86 & new_G4660;
  assign new_G4682 = G109 & new_G4660;
  assign new_G4684 = G110 & new_G4660;
  assign new_G579 = new_G577 & new_G581;
  assign new_G629 = new_G616 & new_G581;
  assign new_G633 = new_G618 & new_G581;
  assign new_G637 = new_G620 & new_G581;
  assign new_G641 = new_G622 & new_G581;
  assign new_G645 = new_G624 & new_G601;
  assign new_G711 = new_G692 & new_G650;
  assign new_G715 = new_G694 & new_G650;
  assign new_G719 = new_G696 & new_G650;
  assign new_G723 = new_G698 & new_G650;
  assign new_G727 = new_G700 & new_G650;
  assign new_G731 = new_G702 & new_G671;
  assign new_G737 = new_G704 & new_G671;
  assign new_G745 = new_G706 & new_G671;
  assign new_G751 = new_G708 & new_G671;
  assign new_G757 = new_G710 & new_G671;
  assign new_G887 = ~new_G885 | ~new_G886;
  assign new_G1019 = ~new_G1017 | ~new_G1018;
  assign new_G5245 = ~new_G5239;
  assign new_G1383 = new_G1365 | new_G1366;
  assign new_G1387 = new_G1367 | new_G1368;
  assign new_G1391 = new_G1369 | new_G1370;
  assign new_G1395 = new_G1371 | new_G1372;
  assign new_G1399 = new_G1375 | new_G1376;
  assign new_G1406 = new_G1377 | new_G1378;
  assign new_G1412 = new_G1379 | new_G1380;
  assign new_G1418 = new_G1381 | new_G1382;
  assign new_G2305 = new_G2287 | new_G2288;
  assign new_G2308 = new_G2289 | new_G2290;
  assign new_G2312 = new_G2291 | new_G2292;
  assign new_G2316 = new_G2293 | new_G2294;
  assign new_G2933 = new_G2920 & new_G2886;
  assign new_G2938 = new_G2922 & new_G2886;
  assign new_G2942 = new_G2924 & new_G2886;
  assign new_G2946 = new_G2926 & new_G2886;
  assign new_G2950 = new_G2928 & new_G2905;
  assign new_G3170 = ~new_G3168 | ~new_G3169;
  assign new_G3210 = ~new_G6554 | ~new_G6557;
  assign new_G3667 = new_G3650 | new_G3651;
  assign new_G3670 = new_G3652 | new_G3653;
  assign new_G3673 = new_G3654 | new_G3655;
  assign new_G3676 = new_G3656 | new_G3657;
  assign new_G3679 = new_G3658 | new_G3659;
  assign new_G3682 = new_G3665 | new_G3635;
  assign new_G3686 = new_G3666 | new_G3635;
  assign new_G3801 = new_G3781 | new_G3782;
  assign new_G3804 = new_G3783 | new_G3784;
  assign new_G3807 = new_G3785 | new_G3786;
  assign new_G3810 = new_G3787 | new_G3788;
  assign new_G3813 = new_G3789 | new_G3790;
  assign new_G4525 = new_G2918 & new_G2886;
  assign new_G4686 = new_G4668 | new_G4669;
  assign new_G4689 = new_G4670 | new_G4671;
  assign new_G4692 = new_G4672 | new_G4673;
  assign new_G4695 = new_G4674 | new_G4675;
  assign new_G4698 = new_G4676 | new_G4677;
  assign new_G4701 = new_G4678 | new_G4679;
  assign new_G4704 = new_G4680 | new_G4681;
  assign new_G4707 = new_G4682 | new_G4683;
  assign new_G4710 = new_G4684 | new_G4685;
  assign new_G4976 = ~new_G4970;
  assign new_G5271 = new_G2932 & new_G2905;
  assign new_G5274 = new_G2930 & new_G2905;
  assign new_G5305 = new_G628 & new_G601;
  assign new_G5308 = new_G626 & new_G601;
  assign new_G5318 = new_G1373 | new_G1374;
  assign new_G6690 = new_G3648 | new_G3649;
  assign new_G6711 = new_G3662 | new_G3663;
  assign new_G6714 = new_G3660 | new_G3661;
  assign new_G7252 = new_G2285 | new_G2286;
  assign new_G7296 = new_G1363 | new_G1364;
  assign new_G7466 = new_G4666 | new_G4667;
  assign new_G907 = new_G765 & new_G784;
  assign new_G913 = new_G765 & new_G784;
  assign new_G915 = new_G765 & new_G784;
  assign new_G916 = new_G765 & new_G784;
  assign new_G1116 = new_G1007 & new_G1014;
  assign new_G2045 = G204 & new_G2026;
  assign new_G2047 = G203 & new_G2026;
  assign new_G2049 = G202 & new_G2026;
  assign new_G2051 = G201 & new_G2026;
  assign new_G2053 = G200 & new_G2026;
  assign new_G2055 = G235 & new_G2039;
  assign new_G2057 = G234 & new_G2039;
  assign new_G2059 = G233 & new_G2039;
  assign new_G2061 = G232 & new_G2039;
  assign new_G2063 = G231 & new_G2039;
  assign new_G2143 = G197 & new_G2124;
  assign new_G2145 = G187 & new_G2124;
  assign new_G2147 = G196 & new_G2124;
  assign new_G2149 = G195 & new_G2124;
  assign new_G2151 = G194 & new_G2124;
  assign new_G2153 = G227 & new_G2137;
  assign new_G2155 = G217 & new_G2137;
  assign new_G2157 = G226 & new_G2137;
  assign new_G2159 = G225 & new_G2137;
  assign new_G2161 = G224 & new_G2137;
  assign new_G2295 = G239 & new_G2279;
  assign new_G2297 = G229 & new_G2279;
  assign new_G2299 = G238 & new_G2279;
  assign new_G2301 = G237 & new_G2279;
  assign new_G2303 = G236 & new_G2279;
  assign new_G3212 = ~new_G3210 | ~new_G3211;
  assign new_G3791 = G223 & new_G3775;
  assign new_G3793 = G222 & new_G3775;
  assign new_G3795 = G221 & new_G3775;
  assign new_G3797 = G220 & new_G3775;
  assign new_G3799 = G219 & new_G3775;
  assign new_G4122 = new_G4121 & new_G4101;
  assign new_G4125 = new_G4396 & new_G4101;
  assign new_G4128 = new_G4402 & new_G4101;
  assign new_G4131 = new_G4407 & new_G4101;
  assign new_G4134 = new_G4412 & new_G4101;
  assign new_G4137 = new_G4417 & new_G4114;
  assign new_G4140 = new_G4422 & new_G4114;
  assign new_G4143 = new_G4429 & new_G4114;
  assign new_G4146 = new_G4434 & new_G4114;
  assign new_G4149 = new_G4439 & new_G4114;
  assign new_G4470 = new_G3700 & new_G4451;
  assign new_G4472 = new_G3703 & new_G4451;
  assign new_G4474 = new_G3707 & new_G4451;
  assign new_G4476 = new_G3713 & new_G4451;
  assign new_G4478 = new_G3719 & new_G4451;
  assign new_G4480 = new_G3725 & new_G4464;
  assign new_G4482 = new_G3731 & new_G4464;
  assign new_G4484 = new_G3739 & new_G4464;
  assign new_G4486 = new_G3745 & new_G4464;
  assign new_G4488 = new_G3751 & new_G4464;
  assign new_G4962 = new_G765;
  assign new_G5003 = new_G765;
  assign new_G5234 = new_G1007;
  assign new_G5242 = new_G1007;
  assign new_G5250 = ~new_G4525;
  assign new_G5284 = ~new_G579;
  assign new_G802 = new_G1488 & new_G2950;
  assign new_G821 = new_G1482 & new_G2946;
  assign new_G845 = new_G1477 & new_G2942;
  assign new_G868 = new_G1471 & new_G2938;
  assign new_G877 = new_G1464 & new_G2933;
  assign new_G902 = new_G887 & new_G765;
  assign new_G908 = new_G777 | new_G907;
  assign new_G914 = new_G887 & new_G765;
  assign new_G917 = new_G777 | new_G916;
  assign new_G953 = new_G887 & new_G765;
  assign new_G1023 = ~new_G1019;
  assign new_G1035 = new_G1488 & new_G2950;
  assign new_G1050 = new_G1482 & new_G2946;
  assign new_G1068 = new_G1477 & new_G2942;
  assign new_G1086 = new_G1471 & new_G2938;
  assign new_G1102 = new_G1464 & new_G2933;
  assign new_G1108 = new_G1019 & new_G1007;
  assign new_G1117 = new_G1115 | new_G1116;
  assign new_G5322 = ~new_G5318;
  assign new_G1553 = new_G1192 & new_G757;
  assign new_G1567 = new_G1186 & new_G751;
  assign new_G1584 = new_G2249 & new_G745;
  assign new_G1590 = new_G2241 & new_G737;
  assign new_G1606 = new_G1178 & new_G731;
  assign new_G1624 = new_G2232 & new_G1418;
  assign new_G1647 = new_G2226 & new_G1412;
  assign new_G1669 = new_G2220 & new_G1406;
  assign new_G1677 = new_G2213 & new_G1399;
  assign new_G1802 = new_G1192 & new_G757;
  assign new_G1816 = new_G1186 & new_G751;
  assign new_G1834 = new_G2249 & new_G745;
  assign new_G1841 = new_G737 & new_G2241;
  assign new_G1866 = new_G1178 & new_G731;
  assign new_G1880 = new_G2232 & new_G1418;
  assign new_G1897 = new_G2226 & new_G1412;
  assign new_G1914 = new_G2220 & new_G1406;
  assign new_G1929 = new_G2213 & new_G1399;
  assign new_G2065 = new_G2045 | new_G2046;
  assign new_G2069 = new_G2047 | new_G2048;
  assign new_G2073 = new_G2049 | new_G2050;
  assign new_G2077 = new_G2051 | new_G2052;
  assign new_G2081 = new_G2053 | new_G2054;
  assign new_G2085 = new_G2055 | new_G2056;
  assign new_G2091 = new_G2057 | new_G2058;
  assign new_G2099 = new_G2059 | new_G2060;
  assign new_G2105 = new_G2061 | new_G2062;
  assign new_G2111 = new_G2063 | new_G2064;
  assign new_G2163 = new_G2145 | new_G2146;
  assign new_G2167 = new_G2147 | new_G2148;
  assign new_G2171 = new_G2149 | new_G2150;
  assign new_G2175 = new_G2151 | new_G2152;
  assign new_G2179 = new_G2155 | new_G2156;
  assign new_G2186 = new_G2157 | new_G2158;
  assign new_G2192 = new_G2159 | new_G2160;
  assign new_G2198 = new_G2161 | new_G2162;
  assign new_G2320 = new_G2297 | new_G2298;
  assign new_G2323 = new_G2299 | new_G2300;
  assign new_G2329 = new_G2301 | new_G2302;
  assign new_G2335 = new_G2303 | new_G2304;
  assign new_G2962 = new_G4710 & new_G727;
  assign new_G2970 = new_G4707 & new_G723;
  assign new_G2977 = new_G4704 & new_G719;
  assign new_G2979 = new_G4701 & new_G715;
  assign new_G2989 = new_G4698 & new_G711;
  assign new_G2998 = new_G4695 & new_G1395;
  assign new_G3006 = new_G4692 & new_G1391;
  assign new_G3013 = new_G4689 & new_G1387;
  assign new_G3015 = new_G4686 & new_G1383;
  assign new_G3183 = new_G3679 & new_G645;
  assign new_G3192 = new_G3676 & new_G641;
  assign new_G3200 = new_G3673 & new_G637;
  assign new_G3207 = new_G3670 & new_G633;
  assign new_G3209 = new_G3667 & new_G629;
  assign new_G3216 = new_G3212 & new_G3170;
  assign new_G3222 = new_G3170 & new_G3173;
  assign new_G6694 = ~new_G6690;
  assign new_G3695 = new_G1535 & new_G2305;
  assign new_G3816 = new_G3791 | new_G3792;
  assign new_G3821 = new_G3793 | new_G3794;
  assign new_G3828 = new_G3795 | new_G3796;
  assign new_G3833 = new_G3797 | new_G3798;
  assign new_G3838 = new_G3799 | new_G3800;
  assign new_G4151 = new_G4125 | new_G4126;
  assign new_G4154 = new_G4128 | new_G4129;
  assign new_G4157 = new_G4131 | new_G4132;
  assign new_G4160 = new_G4134 | new_G4135;
  assign new_G4163 = new_G4137 | new_G4138;
  assign new_G4166 = new_G4140 | new_G4141;
  assign new_G4169 = new_G4143 | new_G4144;
  assign new_G4172 = new_G4146 | new_G4147;
  assign new_G4175 = new_G4149 | new_G4150;
  assign new_G7256 = ~new_G7252;
  assign new_G7300 = ~new_G7296;
  assign new_G4490 = new_G4474 | new_G4475;
  assign new_G4493 = new_G4476 | new_G4477;
  assign new_G4496 = new_G4478 | new_G4479;
  assign new_G4499 = new_G4480 | new_G4481;
  assign new_G4502 = new_G4482 | new_G4483;
  assign new_G4505 = new_G4484 | new_G4485;
  assign new_G4508 = new_G4486 | new_G4487;
  assign new_G4511 = new_G4488 | new_G4489;
  assign new_G7470 = ~new_G7466;
  assign new_G4884 = new_G2950;
  assign new_G4892 = new_G2946;
  assign new_G4900 = new_G2942;
  assign new_G4908 = new_G2938;
  assign new_G4924 = new_G2933;
  assign new_G4952 = new_G887;
  assign new_G4983 = ~new_G777 & ~new_G915;
  assign new_G4993 = new_G887;
  assign new_G5011 = ~new_G1464 & ~new_G2933;
  assign new_G5194 = new_G2950;
  assign new_G5202 = new_G2946;
  assign new_G5210 = new_G2942;
  assign new_G5218 = new_G2938;
  assign new_G5226 = new_G2933;
  assign new_G5247 = new_G2933;
  assign new_G5255 = new_G2942;
  assign new_G5258 = new_G2938;
  assign new_G5263 = new_G2950;
  assign new_G5266 = new_G2946;
  assign new_G5277 = ~new_G5271;
  assign new_G5278 = ~new_G5274;
  assign new_G5281 = new_G629;
  assign new_G5289 = new_G637;
  assign new_G5292 = new_G633;
  assign new_G5297 = new_G645;
  assign new_G5300 = new_G641;
  assign new_G5311 = ~new_G5305;
  assign new_G5312 = ~new_G5308;
  assign new_G5315 = new_G1399;
  assign new_G5323 = new_G1412;
  assign new_G5326 = new_G1406;
  assign new_G5331 = new_G731;
  assign new_G5334 = new_G1418;
  assign new_G5339 = new_G745;
  assign new_G5342 = new_G737;
  assign new_G5349 = new_G757;
  assign new_G5352 = new_G751;
  assign new_G5396 = new_G757;
  assign new_G5404 = new_G751;
  assign new_G5412 = new_G745;
  assign new_G5420 = new_G731;
  assign new_G5428 = new_G1418;
  assign new_G5436 = new_G1412;
  assign new_G5444 = new_G1406;
  assign new_G5452 = new_G737;
  assign new_G5460 = new_G1399;
  assign new_G5465 = ~new_G2241 & ~new_G737;
  assign new_G5581 = ~new_G2213 & ~new_G1399;
  assign new_G5748 = new_G757;
  assign new_G5756 = new_G751;
  assign new_G5764 = new_G745;
  assign new_G5772 = new_G737;
  assign new_G5780 = new_G731;
  assign new_G5788 = new_G1418;
  assign new_G5796 = new_G1412;
  assign new_G5804 = new_G1406;
  assign new_G5812 = new_G1399;
  assign new_G5849 = ~new_G737 & ~new_G2241;
  assign new_G5929 = new_G3682;
  assign new_G6049 = new_G3682;
  assign new_G6367 = new_G4710;
  assign new_G6370 = new_G727;
  assign new_G6375 = new_G4707;
  assign new_G6378 = new_G723;
  assign new_G6383 = new_G4704;
  assign new_G6386 = new_G719;
  assign new_G6391 = new_G4698;
  assign new_G6394 = new_G711;
  assign new_G6399 = new_G4695;
  assign new_G6402 = new_G1395;
  assign new_G6407 = new_G4692;
  assign new_G6410 = new_G1391;
  assign new_G6415 = new_G4689;
  assign new_G6418 = new_G1387;
  assign new_G6423 = new_G4701;
  assign new_G6426 = new_G715;
  assign new_G6431 = new_G4686;
  assign new_G6434 = new_G1383;
  assign new_G6442 = new_G3813;
  assign new_G6450 = new_G3810;
  assign new_G6458 = new_G3807;
  assign new_G6466 = new_G3801;
  assign new_G6498 = new_G3804;
  assign new_G6519 = new_G3679;
  assign new_G6522 = new_G645;
  assign new_G6527 = new_G3676;
  assign new_G6530 = new_G641;
  assign new_G6535 = new_G3673;
  assign new_G6538 = new_G637;
  assign new_G6543 = new_G3670;
  assign new_G6546 = new_G633;
  assign new_G6559 = new_G3667;
  assign new_G6562 = new_G629;
  assign new_G6687 = new_G3667;
  assign new_G6695 = new_G3673;
  assign new_G6698 = new_G3670;
  assign new_G6703 = new_G3679;
  assign new_G6706 = new_G3676;
  assign new_G6717 = ~new_G6711;
  assign new_G6718 = ~new_G6714;
  assign new_G6724 = new_G2153 | new_G2154;
  assign new_G6768 = new_G2295 | new_G2296;
  assign new_G7208 = new_G2143 | new_G2144;
  assign new_G7221 = new_G3801;
  assign new_G7229 = new_G3807;
  assign new_G7232 = new_G3804;
  assign new_G7239 = new_G3813;
  assign new_G7242 = new_G3810;
  assign new_G7249 = new_G2305;
  assign new_G7257 = new_G2312;
  assign new_G7260 = new_G2308;
  assign new_G7268 = new_G2316;
  assign new_G7293 = new_G1383;
  assign new_G7301 = new_G1391;
  assign new_G7304 = new_G1387;
  assign new_G7309 = new_G711;
  assign new_G7312 = new_G1395;
  assign new_G7317 = new_G719;
  assign new_G7320 = new_G715;
  assign new_G7327 = new_G727;
  assign new_G7330 = new_G723;
  assign new_G7396 = new_G2316;
  assign new_G7404 = new_G2312;
  assign new_G7412 = new_G2308;
  assign new_G7425 = new_G3686;
  assign new_G7463 = new_G4686;
  assign new_G7471 = new_G4692;
  assign new_G7474 = new_G4689;
  assign new_G7479 = new_G4698;
  assign new_G7482 = new_G4695;
  assign new_G7487 = new_G4704;
  assign new_G7490 = new_G4701;
  assign new_G7497 = new_G4710;
  assign new_G7500 = new_G4707;
  assign new_G7507 = new_G4472 | new_G4473;
  assign new_G7510 = new_G4470 | new_G4471;
  assign new_G7554 = new_G4122 | new_G4123;
  assign new_G1152 = ~new_G5234 | ~new_G5237;
  assign new_G5238 = ~new_G5234;
  assign new_G1156 = ~new_G5242 | ~new_G5245;
  assign new_G5246 = ~new_G5242;
  assign new_G5254 = ~new_G5250;
  assign new_G5288 = ~new_G5284;
  assign new_G3223 = new_G3221 | new_G3222;
  assign new_G4942 = new_G914 | new_G777 | new_G913;
  assign new_G4966 = ~new_G4962;
  assign new_G5007 = ~new_G5003;
  assign new_G5279 = ~new_G5274 | ~new_G5277;
  assign new_G5280 = ~new_G5271 | ~new_G5278;
  assign new_G5313 = ~new_G5308 | ~new_G5311;
  assign new_G5314 = ~new_G5305 | ~new_G5312;
  assign new_G6719 = ~new_G6714 | ~new_G6717;
  assign new_G6720 = ~new_G6711 | ~new_G6718;
  assign new_G790 = ~new_G4884 | ~new_G4887;
  assign new_G4888 = ~new_G4884;
  assign new_G803 = ~new_G4892 | ~new_G4895;
  assign new_G4896 = ~new_G4892;
  assign new_G825 = ~new_G4900 | ~new_G4903;
  assign new_G4904 = ~new_G4900;
  assign new_G851 = ~new_G4908 | ~new_G4911;
  assign new_G4912 = ~new_G4908;
  assign new_G893 = ~new_G4924 | ~new_G4927;
  assign new_G4928 = ~new_G4924;
  assign new_G906 = ~new_G902;
  assign new_G912 = ~new_G908;
  assign new_G1024 = ~new_G5194 | ~new_G5197;
  assign new_G5198 = ~new_G5194;
  assign new_G1036 = ~new_G5202 | ~new_G5205;
  assign new_G5206 = ~new_G5202;
  assign new_G1053 = ~new_G5210 | ~new_G5213;
  assign new_G5214 = ~new_G5210;
  assign new_G1072 = ~new_G5218 | ~new_G5221;
  assign new_G5222 = ~new_G5218;
  assign new_G1091 = ~new_G5226 | ~new_G5229;
  assign new_G5230 = ~new_G5226;
  assign new_G1112 = ~new_G1108;
  assign new_G1121 = ~new_G1117;
  assign new_G1153 = ~new_G5231 | ~new_G5238;
  assign new_G1157 = ~new_G5239 | ~new_G5246;
  assign new_G5253 = ~new_G5247;
  assign new_G1216 = ~new_G5247 | ~new_G5254;
  assign new_G5261 = ~new_G5255;
  assign new_G5262 = ~new_G5258;
  assign new_G5269 = ~new_G5263;
  assign new_G5270 = ~new_G5266;
  assign new_G5287 = ~new_G5281;
  assign new_G1239 = ~new_G5281 | ~new_G5288;
  assign new_G5295 = ~new_G5289;
  assign new_G5296 = ~new_G5292;
  assign new_G5303 = ~new_G5297;
  assign new_G5304 = ~new_G5300;
  assign new_G5321 = ~new_G5315;
  assign new_G1262 = ~new_G5315 | ~new_G5322;
  assign new_G5329 = ~new_G5323;
  assign new_G5330 = ~new_G5326;
  assign new_G5337 = ~new_G5331;
  assign new_G5338 = ~new_G5334;
  assign new_G1544 = ~new_G5396 | ~new_G5399;
  assign new_G5400 = ~new_G5396;
  assign new_G1554 = ~new_G5404 | ~new_G5407;
  assign new_G5408 = ~new_G5404;
  assign new_G1571 = ~new_G5412 | ~new_G5415;
  assign new_G5416 = ~new_G5412;
  assign new_G1596 = ~new_G5420 | ~new_G5423;
  assign new_G5424 = ~new_G5420;
  assign new_G1607 = ~new_G5428 | ~new_G5431;
  assign new_G5432 = ~new_G5428;
  assign new_G1628 = ~new_G5436 | ~new_G5439;
  assign new_G5440 = ~new_G5436;
  assign new_G1653 = ~new_G5444 | ~new_G5447;
  assign new_G5448 = ~new_G5444;
  assign new_G1685 = ~new_G5452 | ~new_G5455;
  assign new_G5456 = ~new_G5452;
  assign new_G1693 = ~new_G5460 | ~new_G5463;
  assign new_G5464 = ~new_G5460;
  assign new_G1793 = ~new_G5748 | ~new_G5751;
  assign new_G5752 = ~new_G5748;
  assign new_G1803 = ~new_G5756 | ~new_G5759;
  assign new_G5760 = ~new_G5756;
  assign new_G1820 = ~new_G5764 | ~new_G5767;
  assign new_G5768 = ~new_G5764;
  assign new_G1848 = ~new_G5772 | ~new_G5775;
  assign new_G5776 = ~new_G5772;
  assign new_G1857 = ~new_G5780 | ~new_G5783;
  assign new_G5784 = ~new_G5780;
  assign new_G1867 = ~new_G5788 | ~new_G5791;
  assign new_G5792 = ~new_G5788;
  assign new_G1883 = ~new_G5796 | ~new_G5799;
  assign new_G5800 = ~new_G5796;
  assign new_G1901 = ~new_G5804 | ~new_G5807;
  assign new_G5808 = ~new_G5804;
  assign new_G1919 = ~new_G5812 | ~new_G5815;
  assign new_G5816 = ~new_G5812;
  assign new_G5855 = ~new_G5849;
  assign new_G2351 = new_G3751 & new_G2111;
  assign new_G2366 = new_G3745 & new_G2105;
  assign new_G2384 = new_G3739 & new_G2099;
  assign new_G2391 = new_G2091 & new_G3731;
  assign new_G2417 = new_G3725 & new_G2085;
  assign new_G2431 = new_G3719 & new_G2335;
  assign new_G2448 = new_G3713 & new_G2329;
  assign new_G2465 = new_G3707 & new_G2323;
  assign new_G5935 = ~new_G5929;
  assign new_G2597 = new_G3751 & new_G2111;
  assign new_G2612 = new_G3745 & new_G2105;
  assign new_G2629 = new_G3739 & new_G2099;
  assign new_G2635 = new_G3731 & new_G2091;
  assign new_G2652 = new_G3725 & new_G2085;
  assign new_G2670 = new_G3719 & new_G2335;
  assign new_G2693 = new_G3713 & new_G2329;
  assign new_G2715 = new_G3707 & new_G2323;
  assign new_G6055 = ~new_G6049;
  assign new_G6373 = ~new_G6367;
  assign new_G6374 = ~new_G6370;
  assign new_G6381 = ~new_G6375;
  assign new_G6382 = ~new_G6378;
  assign new_G6389 = ~new_G6383;
  assign new_G6390 = ~new_G6386;
  assign new_G6397 = ~new_G6391;
  assign new_G6398 = ~new_G6394;
  assign new_G6405 = ~new_G6399;
  assign new_G6406 = ~new_G6402;
  assign new_G6413 = ~new_G6407;
  assign new_G6414 = ~new_G6410;
  assign new_G6421 = ~new_G6415;
  assign new_G6422 = ~new_G6418;
  assign new_G6429 = ~new_G6423;
  assign new_G6430 = ~new_G6426;
  assign new_G6437 = ~new_G6431;
  assign new_G6438 = ~new_G6434;
  assign new_G6446 = ~new_G6442;
  assign new_G3059 = new_G4175 & new_G3813;
  assign new_G6454 = ~new_G6450;
  assign new_G3068 = new_G4172 & new_G3810;
  assign new_G6462 = ~new_G6458;
  assign new_G3076 = new_G4169 & new_G3807;
  assign new_G3079 = new_G4166 & new_G3804;
  assign new_G6470 = ~new_G6466;
  assign new_G3090 = new_G4163 & new_G3801;
  assign new_G3099 = new_G4160 & new_G2175;
  assign new_G3107 = new_G4157 & new_G2171;
  assign new_G3114 = new_G4154 & new_G2167;
  assign new_G3116 = new_G4151 & new_G2163;
  assign new_G6502 = ~new_G6498;
  assign new_G6525 = ~new_G6519;
  assign new_G6526 = ~new_G6522;
  assign new_G6533 = ~new_G6527;
  assign new_G6534 = ~new_G6530;
  assign new_G6541 = ~new_G6535;
  assign new_G6542 = ~new_G6538;
  assign new_G6549 = ~new_G6543;
  assign new_G6550 = ~new_G6546;
  assign new_G6565 = ~new_G6559;
  assign new_G6566 = ~new_G6562;
  assign new_G3220 = ~new_G3216;
  assign new_G3292 = new_G4439 & new_G3838;
  assign new_G3308 = new_G4434 & new_G3833;
  assign new_G3327 = new_G4429 & new_G3828;
  assign new_G3335 = new_G3821 & new_G4422;
  assign new_G3362 = new_G4417 & new_G3816;
  assign new_G3376 = new_G4412 & new_G2198;
  assign new_G3393 = new_G4407 & new_G2192;
  assign new_G3410 = new_G4402 & new_G2186;
  assign new_G3425 = new_G4396 & new_G2179;
  assign new_G6693 = ~new_G6687;
  assign new_G3503 = ~new_G6687 | ~new_G6694;
  assign new_G6701 = ~new_G6695;
  assign new_G6702 = ~new_G6698;
  assign new_G6709 = ~new_G6703;
  assign new_G6710 = ~new_G6706;
  assign new_G6728 = ~new_G6724;
  assign new_G6772 = ~new_G6768;
  assign new_G3853 = new_G4439 & new_G3838;
  assign new_G3868 = new_G4434 & new_G3833;
  assign new_G3885 = new_G4429 & new_G3828;
  assign new_G3891 = new_G4422 & new_G3821;
  assign new_G3908 = new_G4417 & new_G3816;
  assign new_G3926 = new_G4412 & new_G2198;
  assign new_G3949 = new_G4407 & new_G2192;
  assign new_G3971 = new_G4402 & new_G2186;
  assign new_G3979 = new_G4396 & new_G2179;
  assign new_G7212 = ~new_G7208;
  assign new_G7227 = ~new_G7221;
  assign new_G7255 = ~new_G7249;
  assign new_G4202 = ~new_G7249 | ~new_G7256;
  assign new_G7263 = ~new_G7257;
  assign new_G7264 = ~new_G7260;
  assign new_G7272 = ~new_G7268;
  assign new_G7299 = ~new_G7293;
  assign new_G4225 = ~new_G7293 | ~new_G7300;
  assign new_G7307 = ~new_G7301;
  assign new_G7308 = ~new_G7304;
  assign new_G7315 = ~new_G7309;
  assign new_G7316 = ~new_G7312;
  assign new_G4297 = new_G4511 & new_G2081;
  assign new_G4305 = new_G4508 & new_G2077;
  assign new_G4312 = new_G4505 & new_G2073;
  assign new_G4314 = new_G4502 & new_G2069;
  assign new_G4324 = new_G4499 & new_G2065;
  assign new_G7400 = ~new_G7396;
  assign new_G4333 = new_G4496 & new_G2316;
  assign new_G7408 = ~new_G7404;
  assign new_G4341 = new_G4493 & new_G2312;
  assign new_G7416 = ~new_G7412;
  assign new_G4348 = new_G4490 & new_G2308;
  assign new_G4349 = new_G3686 & new_G3695;
  assign new_G7431 = ~new_G7425;
  assign new_G4389 = new_G2320 & new_G1535;
  assign new_G7469 = ~new_G7463;
  assign new_G4530 = ~new_G7463 | ~new_G7470;
  assign new_G7477 = ~new_G7471;
  assign new_G7478 = ~new_G7474;
  assign new_G7485 = ~new_G7479;
  assign new_G7486 = ~new_G7482;
  assign new_G7513 = ~new_G7507;
  assign new_G7514 = ~new_G7510;
  assign new_G7558 = ~new_G7554;
  assign new_G4932 = new_G917 | new_G953;
  assign new_G4956 = ~new_G4952;
  assign new_G4973 = ~new_G917;
  assign new_G4987 = ~new_G4983;
  assign new_G4997 = ~new_G4993;
  assign new_G5017 = ~new_G5011;
  assign new_G5099 = new_G877;
  assign new_G5345 = ~new_G5339;
  assign new_G5346 = ~new_G5342;
  assign new_G5355 = ~new_G5349;
  assign new_G5356 = ~new_G5352;
  assign new_G5372 = ~new_G5279 | ~new_G5280;
  assign new_G5380 = ~new_G5313 | ~new_G5314;
  assign new_G5471 = ~new_G5465;
  assign new_G5523 = new_G1590;
  assign new_G5587 = ~new_G5581;
  assign new_G5669 = new_G1677;
  assign new_G5857 = new_G1841;
  assign new_G5868 = new_G2111;
  assign new_G5876 = new_G2105;
  assign new_G5884 = new_G2099;
  assign new_G5892 = new_G2091;
  assign new_G5900 = new_G2085;
  assign new_G5908 = new_G2335;
  assign new_G5916 = new_G2329;
  assign new_G5924 = new_G2323;
  assign new_G5969 = ~new_G2091 & ~new_G3731;
  assign new_G5988 = new_G2111;
  assign new_G5996 = new_G2105;
  assign new_G6004 = new_G2099;
  assign new_G6012 = new_G2085;
  assign new_G6020 = new_G2335;
  assign new_G6028 = new_G2329;
  assign new_G6036 = new_G2323;
  assign new_G6044 = new_G2091;
  assign new_G6057 = ~new_G3731 & ~new_G2091;
  assign new_G6439 = new_G4175;
  assign new_G6447 = new_G4172;
  assign new_G6455 = new_G4169;
  assign new_G6463 = new_G4163;
  assign new_G6471 = new_G4160;
  assign new_G6474 = new_G2175;
  assign new_G6479 = new_G4157;
  assign new_G6482 = new_G2171;
  assign new_G6487 = new_G4154;
  assign new_G6490 = new_G2167;
  assign new_G6495 = new_G4166;
  assign new_G6503 = new_G4151;
  assign new_G6506 = new_G2163;
  assign new_G6570 = new_G3838;
  assign new_G6578 = new_G3833;
  assign new_G6586 = new_G3828;
  assign new_G6594 = new_G3821;
  assign new_G6602 = new_G3816;
  assign new_G6610 = new_G2198;
  assign new_G6618 = new_G2192;
  assign new_G6626 = new_G2186;
  assign new_G6634 = new_G2179;
  assign new_G6671 = ~new_G3821 & ~new_G4422;
  assign new_G6721 = new_G2179;
  assign new_G6729 = new_G2192;
  assign new_G6732 = new_G2186;
  assign new_G6737 = new_G3816;
  assign new_G6740 = new_G2198;
  assign new_G6745 = new_G3828;
  assign new_G6748 = new_G3821;
  assign new_G6755 = new_G3838;
  assign new_G6758 = new_G3833;
  assign new_G6765 = new_G2320;
  assign new_G6773 = new_G2329;
  assign new_G6776 = new_G2323;
  assign new_G6781 = new_G2085;
  assign new_G6784 = new_G2335;
  assign new_G6789 = new_G2099;
  assign new_G6792 = new_G2091;
  assign new_G6799 = new_G2111;
  assign new_G6802 = new_G2105;
  assign new_G6832 = ~new_G6719 | ~new_G6720;
  assign new_G6856 = new_G3838;
  assign new_G6864 = new_G3833;
  assign new_G6872 = new_G3828;
  assign new_G6880 = new_G3816;
  assign new_G6888 = new_G2198;
  assign new_G6896 = new_G2192;
  assign new_G6904 = new_G2186;
  assign new_G6912 = new_G3821;
  assign new_G6920 = new_G2179;
  assign new_G6925 = ~new_G4422 & ~new_G3821;
  assign new_G7041 = ~new_G4396 & ~new_G2179;
  assign new_G7205 = new_G2163;
  assign new_G7213 = new_G2171;
  assign new_G7216 = new_G2167;
  assign new_G7224 = new_G2175;
  assign new_G7235 = ~new_G7229;
  assign new_G7236 = ~new_G7232;
  assign new_G7245 = ~new_G7239;
  assign new_G7246 = ~new_G7242;
  assign new_G7265 = new_G2065;
  assign new_G7273 = new_G2073;
  assign new_G7276 = new_G2069;
  assign new_G7283 = new_G2081;
  assign new_G7286 = new_G2077;
  assign new_G7323 = ~new_G7317;
  assign new_G7324 = ~new_G7320;
  assign new_G7333 = ~new_G7327;
  assign new_G7334 = ~new_G7330;
  assign new_G7361 = new_G4511;
  assign new_G7364 = new_G2081;
  assign new_G7369 = new_G4508;
  assign new_G7372 = new_G2077;
  assign new_G7377 = new_G4505;
  assign new_G7380 = new_G2073;
  assign new_G7385 = new_G4499;
  assign new_G7388 = new_G2065;
  assign new_G7393 = new_G4496;
  assign new_G7401 = new_G4493;
  assign new_G7409 = new_G4490;
  assign new_G7417 = new_G4502;
  assign new_G7420 = new_G2069;
  assign new_G7428 = new_G3695;
  assign new_G7493 = ~new_G7487;
  assign new_G7494 = ~new_G7490;
  assign new_G7503 = ~new_G7497;
  assign new_G7504 = ~new_G7500;
  assign new_G7515 = new_G4493;
  assign new_G7518 = new_G4490;
  assign new_G7523 = new_G4499;
  assign new_G7526 = new_G4496;
  assign new_G7531 = new_G4505;
  assign new_G7534 = new_G4502;
  assign new_G7541 = new_G4511;
  assign new_G7544 = new_G4508;
  assign new_G7551 = new_G4151;
  assign new_G7559 = new_G4157;
  assign new_G7562 = new_G4154;
  assign new_G7567 = new_G4163;
  assign new_G7570 = new_G4160;
  assign new_G7575 = new_G4169;
  assign new_G7578 = new_G4166;
  assign new_G7585 = new_G4175;
  assign new_G7588 = new_G4172;
  assign new_G1176 = ~new_G1121 | ~new_G1112;
  assign new_G957 = ~new_G912 | ~new_G906;
  assign new_G791 = ~new_G4881 | ~new_G4888;
  assign new_G804 = ~new_G4889 | ~new_G4896;
  assign new_G826 = ~new_G4897 | ~new_G4904;
  assign new_G852 = ~new_G4905 | ~new_G4912;
  assign new_G894 = ~new_G4921 | ~new_G4928;
  assign new_G1025 = ~new_G5191 | ~new_G5198;
  assign new_G1037 = ~new_G5199 | ~new_G5206;
  assign new_G1054 = ~new_G5207 | ~new_G5214;
  assign new_G1073 = ~new_G5215 | ~new_G5222;
  assign new_G1092 = ~new_G5223 | ~new_G5230;
  assign new_G1154 = ~new_G1152 | ~new_G1153;
  assign new_G1158 = ~new_G1156 | ~new_G1157;
  assign new_G1215 = ~new_G5250 | ~new_G5253;
  assign new_G1224 = ~new_G5258 | ~new_G5261;
  assign new_G1225 = ~new_G5255 | ~new_G5262;
  assign new_G1233 = ~new_G5266 | ~new_G5269;
  assign new_G1234 = ~new_G5263 | ~new_G5270;
  assign new_G1238 = ~new_G5284 | ~new_G5287;
  assign new_G1247 = ~new_G5292 | ~new_G5295;
  assign new_G1248 = ~new_G5289 | ~new_G5296;
  assign new_G1256 = ~new_G5300 | ~new_G5303;
  assign new_G1257 = ~new_G5297 | ~new_G5304;
  assign new_G1261 = ~new_G5318 | ~new_G5321;
  assign new_G1270 = ~new_G5326 | ~new_G5329;
  assign new_G1271 = ~new_G5323 | ~new_G5330;
  assign new_G1279 = ~new_G5334 | ~new_G5337;
  assign new_G1280 = ~new_G5331 | ~new_G5338;
  assign new_G1545 = ~new_G5393 | ~new_G5400;
  assign new_G1555 = ~new_G5401 | ~new_G5408;
  assign new_G1572 = ~new_G5409 | ~new_G5416;
  assign new_G1597 = ~new_G5417 | ~new_G5424;
  assign new_G1608 = ~new_G5425 | ~new_G5432;
  assign new_G1629 = ~new_G5433 | ~new_G5440;
  assign new_G1654 = ~new_G5441 | ~new_G5448;
  assign new_G1686 = ~new_G5449 | ~new_G5456;
  assign new_G1694 = ~new_G5457 | ~new_G5464;
  assign new_G1794 = ~new_G5745 | ~new_G5752;
  assign new_G1804 = ~new_G5753 | ~new_G5760;
  assign new_G1821 = ~new_G5761 | ~new_G5768;
  assign new_G1849 = ~new_G5769 | ~new_G5776;
  assign new_G1858 = ~new_G5777 | ~new_G5784;
  assign new_G1868 = ~new_G5785 | ~new_G5792;
  assign new_G1884 = ~new_G5793 | ~new_G5800;
  assign new_G1902 = ~new_G5801 | ~new_G5808;
  assign new_G1920 = ~new_G5809 | ~new_G5816;
  assign new_G2954 = ~new_G6370 | ~new_G6373;
  assign new_G2955 = ~new_G6367 | ~new_G6374;
  assign new_G2963 = ~new_G6378 | ~new_G6381;
  assign new_G2964 = ~new_G6375 | ~new_G6382;
  assign new_G2971 = ~new_G6386 | ~new_G6389;
  assign new_G2972 = ~new_G6383 | ~new_G6390;
  assign new_G2980 = ~new_G6394 | ~new_G6397;
  assign new_G2981 = ~new_G6391 | ~new_G6398;
  assign new_G2990 = ~new_G6402 | ~new_G6405;
  assign new_G2991 = ~new_G6399 | ~new_G6406;
  assign new_G2999 = ~new_G6410 | ~new_G6413;
  assign new_G3000 = ~new_G6407 | ~new_G6414;
  assign new_G3007 = ~new_G6418 | ~new_G6421;
  assign new_G3008 = ~new_G6415 | ~new_G6422;
  assign new_G3016 = ~new_G6426 | ~new_G6429;
  assign new_G3017 = ~new_G6423 | ~new_G6430;
  assign new_G3019 = ~new_G6434 | ~new_G6437;
  assign new_G3020 = ~new_G6431 | ~new_G6438;
  assign new_G3174 = ~new_G6522 | ~new_G6525;
  assign new_G3175 = ~new_G6519 | ~new_G6526;
  assign new_G3184 = ~new_G6530 | ~new_G6533;
  assign new_G3185 = ~new_G6527 | ~new_G6534;
  assign new_G3193 = ~new_G6538 | ~new_G6541;
  assign new_G3194 = ~new_G6535 | ~new_G6542;
  assign new_G3201 = ~new_G6546 | ~new_G6549;
  assign new_G3202 = ~new_G6543 | ~new_G6550;
  assign new_G3213 = ~new_G6562 | ~new_G6565;
  assign new_G3214 = ~new_G6559 | ~new_G6566;
  assign new_G3227 = ~new_G3223;
  assign new_G3502 = ~new_G6690 | ~new_G6693;
  assign new_G3511 = ~new_G6698 | ~new_G6701;
  assign new_G3512 = ~new_G6695 | ~new_G6702;
  assign new_G3520 = ~new_G6706 | ~new_G6709;
  assign new_G3521 = ~new_G6703 | ~new_G6710;
  assign new_G4201 = ~new_G7252 | ~new_G7255;
  assign new_G4210 = ~new_G7260 | ~new_G7263;
  assign new_G4211 = ~new_G7257 | ~new_G7264;
  assign new_G4224 = ~new_G7296 | ~new_G7299;
  assign new_G4233 = ~new_G7304 | ~new_G7307;
  assign new_G4234 = ~new_G7301 | ~new_G7308;
  assign new_G4242 = ~new_G7312 | ~new_G7315;
  assign new_G4243 = ~new_G7309 | ~new_G7316;
  assign new_G4529 = ~new_G7466 | ~new_G7469;
  assign new_G4538 = ~new_G7474 | ~new_G7477;
  assign new_G4539 = ~new_G7471 | ~new_G7478;
  assign new_G4547 = ~new_G7482 | ~new_G7485;
  assign new_G4548 = ~new_G7479 | ~new_G7486;
  assign new_G4552 = ~new_G7510 | ~new_G7513;
  assign new_G4553 = ~new_G7507 | ~new_G7514;
  assign new_G4946 = ~new_G4942;
  assign new_G5347 = ~new_G5342 | ~new_G5345;
  assign new_G5348 = ~new_G5339 | ~new_G5346;
  assign new_G5357 = ~new_G5352 | ~new_G5355;
  assign new_G5358 = ~new_G5349 | ~new_G5356;
  assign new_G7237 = ~new_G7232 | ~new_G7235;
  assign new_G7238 = ~new_G7229 | ~new_G7236;
  assign new_G7247 = ~new_G7242 | ~new_G7245;
  assign new_G7248 = ~new_G7239 | ~new_G7246;
  assign new_G7325 = ~new_G7320 | ~new_G7323;
  assign new_G7326 = ~new_G7317 | ~new_G7324;
  assign new_G7335 = ~new_G7330 | ~new_G7333;
  assign new_G7336 = ~new_G7327 | ~new_G7334;
  assign new_G7495 = ~new_G7490 | ~new_G7493;
  assign new_G7496 = ~new_G7487 | ~new_G7494;
  assign new_G7505 = ~new_G7500 | ~new_G7503;
  assign new_G7506 = ~new_G7497 | ~new_G7504;
  assign new_G3244 = ~new_G3227 | ~new_G3220;
  assign new_G792 = ~new_G790 | ~new_G791;
  assign new_G805 = ~new_G803 | ~new_G804;
  assign new_G827 = ~new_G825 | ~new_G826;
  assign new_G853 = ~new_G851 | ~new_G852;
  assign new_G895 = ~new_G893 | ~new_G894;
  assign new_G1026 = ~new_G1024 | ~new_G1025;
  assign new_G1038 = ~new_G1036 | ~new_G1037;
  assign new_G1055 = ~new_G1053 | ~new_G1054;
  assign new_G1074 = ~new_G1072 | ~new_G1073;
  assign new_G1093 = ~new_G1091 | ~new_G1092;
  assign new_G1155 = ~new_G1154;
  assign new_G1217 = ~new_G1215 | ~new_G1216;
  assign new_G1226 = ~new_G1224 | ~new_G1225;
  assign new_G1235 = ~new_G1233 | ~new_G1234;
  assign new_G1240 = ~new_G1238 | ~new_G1239;
  assign new_G1249 = ~new_G1247 | ~new_G1248;
  assign new_G1258 = ~new_G1256 | ~new_G1257;
  assign new_G1263 = ~new_G1261 | ~new_G1262;
  assign new_G1272 = ~new_G1270 | ~new_G1271;
  assign new_G1281 = ~new_G1279 | ~new_G1280;
  assign new_G5376 = ~new_G5372;
  assign new_G5384 = ~new_G5380;
  assign new_G1546 = ~new_G1544 | ~new_G1545;
  assign new_G1556 = ~new_G1554 | ~new_G1555;
  assign new_G1573 = ~new_G1571 | ~new_G1572;
  assign new_G1598 = ~new_G1596 | ~new_G1597;
  assign new_G1609 = ~new_G1607 | ~new_G1608;
  assign new_G1630 = ~new_G1628 | ~new_G1629;
  assign new_G1655 = ~new_G1653 | ~new_G1654;
  assign new_G1687 = ~new_G1685 | ~new_G1686;
  assign new_G1695 = ~new_G1693 | ~new_G1694;
  assign new_G1795 = ~new_G1793 | ~new_G1794;
  assign new_G1805 = ~new_G1803 | ~new_G1804;
  assign new_G1822 = ~new_G1820 | ~new_G1821;
  assign new_G1850 = ~new_G1848 | ~new_G1849;
  assign new_G1859 = ~new_G1857 | ~new_G1858;
  assign new_G1869 = ~new_G1867 | ~new_G1868;
  assign new_G1885 = ~new_G1883 | ~new_G1884;
  assign new_G1903 = ~new_G1901 | ~new_G1902;
  assign new_G1921 = ~new_G1919 | ~new_G1920;
  assign new_G5863 = ~new_G5857;
  assign new_G2341 = ~new_G5868 | ~new_G5871;
  assign new_G5872 = ~new_G5868;
  assign new_G2352 = ~new_G5876 | ~new_G5879;
  assign new_G5880 = ~new_G5876;
  assign new_G2370 = ~new_G5884 | ~new_G5887;
  assign new_G5888 = ~new_G5884;
  assign new_G2398 = ~new_G5892 | ~new_G5895;
  assign new_G5896 = ~new_G5892;
  assign new_G2407 = ~new_G5900 | ~new_G5903;
  assign new_G5904 = ~new_G5900;
  assign new_G2418 = ~new_G5908 | ~new_G5911;
  assign new_G5912 = ~new_G5908;
  assign new_G2434 = ~new_G5916 | ~new_G5919;
  assign new_G5920 = ~new_G5916;
  assign new_G2452 = ~new_G5924 | ~new_G5927;
  assign new_G5928 = ~new_G5924;
  assign new_G2481 = new_G3682 & new_G4389;
  assign new_G5975 = ~new_G5969;
  assign new_G2587 = ~new_G5988 | ~new_G5991;
  assign new_G5992 = ~new_G5988;
  assign new_G2598 = ~new_G5996 | ~new_G5999;
  assign new_G6000 = ~new_G5996;
  assign new_G2616 = ~new_G6004 | ~new_G6007;
  assign new_G6008 = ~new_G6004;
  assign new_G2641 = ~new_G6012 | ~new_G6015;
  assign new_G6016 = ~new_G6012;
  assign new_G2653 = ~new_G6020 | ~new_G6023;
  assign new_G6024 = ~new_G6020;
  assign new_G2674 = ~new_G6028 | ~new_G6031;
  assign new_G6032 = ~new_G6028;
  assign new_G2699 = ~new_G6036 | ~new_G6039;
  assign new_G6040 = ~new_G6036;
  assign new_G2724 = new_G3682 & new_G4389;
  assign new_G2732 = ~new_G6044 | ~new_G6047;
  assign new_G6048 = ~new_G6044;
  assign new_G2956 = ~new_G2954 | ~new_G2955;
  assign new_G2965 = ~new_G2963 | ~new_G2964;
  assign new_G2973 = ~new_G2971 | ~new_G2972;
  assign new_G2982 = ~new_G2980 | ~new_G2981;
  assign new_G2992 = ~new_G2990 | ~new_G2991;
  assign new_G3001 = ~new_G2999 | ~new_G3000;
  assign new_G3009 = ~new_G3007 | ~new_G3008;
  assign new_G3018 = ~new_G3016 | ~new_G3017;
  assign new_G3021 = ~new_G3019 | ~new_G3020;
  assign new_G6445 = ~new_G6439;
  assign new_G3051 = ~new_G6439 | ~new_G6446;
  assign new_G6453 = ~new_G6447;
  assign new_G3061 = ~new_G6447 | ~new_G6454;
  assign new_G6461 = ~new_G6455;
  assign new_G3070 = ~new_G6455 | ~new_G6462;
  assign new_G6469 = ~new_G6463;
  assign new_G3081 = ~new_G6463 | ~new_G6470;
  assign new_G6477 = ~new_G6471;
  assign new_G6478 = ~new_G6474;
  assign new_G6485 = ~new_G6479;
  assign new_G6486 = ~new_G6482;
  assign new_G6493 = ~new_G6487;
  assign new_G6494 = ~new_G6490;
  assign new_G6501 = ~new_G6495;
  assign new_G3118 = ~new_G6495 | ~new_G6502;
  assign new_G6509 = ~new_G6503;
  assign new_G6510 = ~new_G6506;
  assign new_G3176 = ~new_G3174 | ~new_G3175;
  assign new_G3186 = ~new_G3184 | ~new_G3185;
  assign new_G3195 = ~new_G3193 | ~new_G3194;
  assign new_G3203 = ~new_G3201 | ~new_G3202;
  assign new_G3215 = ~new_G3213 | ~new_G3214;
  assign new_G3281 = ~new_G6570 | ~new_G6573;
  assign new_G6574 = ~new_G6570;
  assign new_G3293 = ~new_G6578 | ~new_G6581;
  assign new_G6582 = ~new_G6578;
  assign new_G3312 = ~new_G6586 | ~new_G6589;
  assign new_G6590 = ~new_G6586;
  assign new_G3342 = ~new_G6594 | ~new_G6597;
  assign new_G6598 = ~new_G6594;
  assign new_G3351 = ~new_G6602 | ~new_G6605;
  assign new_G6606 = ~new_G6602;
  assign new_G3363 = ~new_G6610 | ~new_G6613;
  assign new_G6614 = ~new_G6610;
  assign new_G3379 = ~new_G6618 | ~new_G6621;
  assign new_G6622 = ~new_G6618;
  assign new_G3397 = ~new_G6626 | ~new_G6629;
  assign new_G6630 = ~new_G6626;
  assign new_G3415 = ~new_G6634 | ~new_G6637;
  assign new_G6638 = ~new_G6634;
  assign new_G6677 = ~new_G6671;
  assign new_G3504 = ~new_G3502 | ~new_G3503;
  assign new_G3513 = ~new_G3511 | ~new_G3512;
  assign new_G3522 = ~new_G3520 | ~new_G3521;
  assign new_G6727 = ~new_G6721;
  assign new_G3526 = ~new_G6721 | ~new_G6728;
  assign new_G6735 = ~new_G6729;
  assign new_G6736 = ~new_G6732;
  assign new_G6743 = ~new_G6737;
  assign new_G6744 = ~new_G6740;
  assign new_G6771 = ~new_G6765;
  assign new_G3549 = ~new_G6765 | ~new_G6772;
  assign new_G6779 = ~new_G6773;
  assign new_G6780 = ~new_G6776;
  assign new_G6787 = ~new_G6781;
  assign new_G6788 = ~new_G6784;
  assign new_G6836 = ~new_G6832;
  assign new_G3843 = ~new_G6856 | ~new_G6859;
  assign new_G6860 = ~new_G6856;
  assign new_G3854 = ~new_G6864 | ~new_G6867;
  assign new_G6868 = ~new_G6864;
  assign new_G3872 = ~new_G6872 | ~new_G6875;
  assign new_G6876 = ~new_G6872;
  assign new_G3897 = ~new_G6880 | ~new_G6883;
  assign new_G6884 = ~new_G6880;
  assign new_G3909 = ~new_G6888 | ~new_G6891;
  assign new_G6892 = ~new_G6888;
  assign new_G3930 = ~new_G6896 | ~new_G6899;
  assign new_G6900 = ~new_G6896;
  assign new_G3955 = ~new_G6904 | ~new_G6907;
  assign new_G6908 = ~new_G6904;
  assign new_G3987 = ~new_G6912 | ~new_G6915;
  assign new_G6916 = ~new_G6912;
  assign new_G3995 = ~new_G6920 | ~new_G6923;
  assign new_G6924 = ~new_G6920;
  assign new_G7211 = ~new_G7205;
  assign new_G4179 = ~new_G7205 | ~new_G7212;
  assign new_G7219 = ~new_G7213;
  assign new_G7220 = ~new_G7216;
  assign new_G4196 = ~new_G7224 | ~new_G7227;
  assign new_G7228 = ~new_G7224;
  assign new_G4203 = ~new_G4201 | ~new_G4202;
  assign new_G4212 = ~new_G4210 | ~new_G4211;
  assign new_G7271 = ~new_G7265;
  assign new_G4220 = ~new_G7265 | ~new_G7272;
  assign new_G4226 = ~new_G4224 | ~new_G4225;
  assign new_G4235 = ~new_G4233 | ~new_G4234;
  assign new_G4244 = ~new_G4242 | ~new_G4243;
  assign new_G7367 = ~new_G7361;
  assign new_G7368 = ~new_G7364;
  assign new_G7375 = ~new_G7369;
  assign new_G7376 = ~new_G7372;
  assign new_G7383 = ~new_G7377;
  assign new_G7384 = ~new_G7380;
  assign new_G7391 = ~new_G7385;
  assign new_G7392 = ~new_G7388;
  assign new_G7399 = ~new_G7393;
  assign new_G4326 = ~new_G7393 | ~new_G7400;
  assign new_G7407 = ~new_G7401;
  assign new_G4335 = ~new_G7401 | ~new_G7408;
  assign new_G7415 = ~new_G7409;
  assign new_G4343 = ~new_G7409 | ~new_G7416;
  assign new_G7423 = ~new_G7417;
  assign new_G7424 = ~new_G7420;
  assign new_G4353 = ~new_G7428 | ~new_G7431;
  assign new_G7432 = ~new_G7428;
  assign new_G4531 = ~new_G4529 | ~new_G4530;
  assign new_G4540 = ~new_G4538 | ~new_G4539;
  assign new_G4549 = ~new_G4547 | ~new_G4548;
  assign new_G4554 = ~new_G4552 | ~new_G4553;
  assign new_G7521 = ~new_G7515;
  assign new_G7522 = ~new_G7518;
  assign new_G7529 = ~new_G7523;
  assign new_G7530 = ~new_G7526;
  assign new_G7557 = ~new_G7551;
  assign new_G4576 = ~new_G7551 | ~new_G7558;
  assign new_G7565 = ~new_G7559;
  assign new_G7566 = ~new_G7562;
  assign new_G7573 = ~new_G7567;
  assign new_G7574 = ~new_G7570;
  assign new_G4936 = ~new_G4932;
  assign new_G4937 = ~new_G4932 | ~new_G4935;
  assign new_G4977 = ~new_G4973;
  assign new_G4978 = ~new_G4973 | ~new_G4976;
  assign new_G5105 = ~new_G5099;
  assign new_G5359 = ~new_G5357 | ~new_G5358;
  assign new_G5362 = ~new_G5347 | ~new_G5348;
  assign new_G5529 = ~new_G5523;
  assign new_G5675 = ~new_G5669;
  assign new_G5932 = new_G4389;
  assign new_G5977 = new_G2391;
  assign new_G6052 = new_G4389;
  assign new_G6063 = ~new_G6057;
  assign new_G6115 = new_G2635;
  assign new_G6173 = ~new_G3682 & ~new_G4389;
  assign new_G6679 = new_G3335;
  assign new_G6751 = ~new_G6745;
  assign new_G6752 = ~new_G6748;
  assign new_G6761 = ~new_G6755;
  assign new_G6762 = ~new_G6758;
  assign new_G6795 = ~new_G6789;
  assign new_G6796 = ~new_G6792;
  assign new_G6805 = ~new_G6799;
  assign new_G6806 = ~new_G6802;
  assign new_G6931 = ~new_G6925;
  assign new_G6983 = new_G3891;
  assign new_G7047 = ~new_G7041;
  assign new_G7129 = new_G3979;
  assign new_G7279 = ~new_G7273;
  assign new_G7280 = ~new_G7276;
  assign new_G7289 = ~new_G7283;
  assign new_G7290 = ~new_G7286;
  assign new_G7337 = ~new_G7247 | ~new_G7248;
  assign new_G7340 = ~new_G7237 | ~new_G7238;
  assign new_G7353 = ~new_G7335 | ~new_G7336;
  assign new_G7356 = ~new_G7325 | ~new_G7326;
  assign new_G7537 = ~new_G7531;
  assign new_G7538 = ~new_G7534;
  assign new_G7547 = ~new_G7541;
  assign new_G7548 = ~new_G7544;
  assign new_G7581 = ~new_G7575;
  assign new_G7582 = ~new_G7578;
  assign new_G7591 = ~new_G7585;
  assign new_G7592 = ~new_G7588;
  assign new_G7595 = ~new_G7505 | ~new_G7506;
  assign new_G7598 = ~new_G7495 | ~new_G7496;
  assign new_G2342 = ~new_G5865 | ~new_G5872;
  assign new_G2353 = ~new_G5873 | ~new_G5880;
  assign new_G2371 = ~new_G5881 | ~new_G5888;
  assign new_G2399 = ~new_G5889 | ~new_G5896;
  assign new_G2408 = ~new_G5897 | ~new_G5904;
  assign new_G2419 = ~new_G5905 | ~new_G5912;
  assign new_G2435 = ~new_G5913 | ~new_G5920;
  assign new_G2453 = ~new_G5921 | ~new_G5928;
  assign new_G2588 = ~new_G5985 | ~new_G5992;
  assign new_G2599 = ~new_G5993 | ~new_G6000;
  assign new_G2617 = ~new_G6001 | ~new_G6008;
  assign new_G2642 = ~new_G6009 | ~new_G6016;
  assign new_G2654 = ~new_G6017 | ~new_G6024;
  assign new_G2675 = ~new_G6025 | ~new_G6032;
  assign new_G2700 = ~new_G6033 | ~new_G6040;
  assign new_G2733 = ~new_G6041 | ~new_G6048;
  assign new_G3050 = ~new_G6442 | ~new_G6445;
  assign new_G3060 = ~new_G6450 | ~new_G6453;
  assign new_G3069 = ~new_G6458 | ~new_G6461;
  assign new_G3080 = ~new_G6466 | ~new_G6469;
  assign new_G3091 = ~new_G6474 | ~new_G6477;
  assign new_G3092 = ~new_G6471 | ~new_G6478;
  assign new_G3100 = ~new_G6482 | ~new_G6485;
  assign new_G3101 = ~new_G6479 | ~new_G6486;
  assign new_G3108 = ~new_G6490 | ~new_G6493;
  assign new_G3109 = ~new_G6487 | ~new_G6494;
  assign new_G3117 = ~new_G6498 | ~new_G6501;
  assign new_G3120 = ~new_G6506 | ~new_G6509;
  assign new_G3121 = ~new_G6503 | ~new_G6510;
  assign new_G3282 = ~new_G6567 | ~new_G6574;
  assign new_G3294 = ~new_G6575 | ~new_G6582;
  assign new_G3313 = ~new_G6583 | ~new_G6590;
  assign new_G3343 = ~new_G6591 | ~new_G6598;
  assign new_G3352 = ~new_G6599 | ~new_G6606;
  assign new_G3364 = ~new_G6607 | ~new_G6614;
  assign new_G3380 = ~new_G6615 | ~new_G6622;
  assign new_G3398 = ~new_G6623 | ~new_G6630;
  assign new_G3416 = ~new_G6631 | ~new_G6638;
  assign new_G3525 = ~new_G6724 | ~new_G6727;
  assign new_G3534 = ~new_G6732 | ~new_G6735;
  assign new_G3535 = ~new_G6729 | ~new_G6736;
  assign new_G3543 = ~new_G6740 | ~new_G6743;
  assign new_G3544 = ~new_G6737 | ~new_G6744;
  assign new_G3548 = ~new_G6768 | ~new_G6771;
  assign new_G3557 = ~new_G6776 | ~new_G6779;
  assign new_G3558 = ~new_G6773 | ~new_G6780;
  assign new_G3566 = ~new_G6784 | ~new_G6787;
  assign new_G3567 = ~new_G6781 | ~new_G6788;
  assign new_G3844 = ~new_G6853 | ~new_G6860;
  assign new_G3855 = ~new_G6861 | ~new_G6868;
  assign new_G3873 = ~new_G6869 | ~new_G6876;
  assign new_G3898 = ~new_G6877 | ~new_G6884;
  assign new_G3910 = ~new_G6885 | ~new_G6892;
  assign new_G3931 = ~new_G6893 | ~new_G6900;
  assign new_G3956 = ~new_G6901 | ~new_G6908;
  assign new_G3988 = ~new_G6909 | ~new_G6916;
  assign new_G3996 = ~new_G6917 | ~new_G6924;
  assign new_G4178 = ~new_G7208 | ~new_G7211;
  assign new_G4187 = ~new_G7216 | ~new_G7219;
  assign new_G4188 = ~new_G7213 | ~new_G7220;
  assign new_G4197 = ~new_G7221 | ~new_G7228;
  assign new_G4219 = ~new_G7268 | ~new_G7271;
  assign new_G4289 = ~new_G7364 | ~new_G7367;
  assign new_G4290 = ~new_G7361 | ~new_G7368;
  assign new_G4298 = ~new_G7372 | ~new_G7375;
  assign new_G4299 = ~new_G7369 | ~new_G7376;
  assign new_G4306 = ~new_G7380 | ~new_G7383;
  assign new_G4307 = ~new_G7377 | ~new_G7384;
  assign new_G4315 = ~new_G7388 | ~new_G7391;
  assign new_G4316 = ~new_G7385 | ~new_G7392;
  assign new_G4325 = ~new_G7396 | ~new_G7399;
  assign new_G4334 = ~new_G7404 | ~new_G7407;
  assign new_G4342 = ~new_G7412 | ~new_G7415;
  assign new_G4350 = ~new_G7420 | ~new_G7423;
  assign new_G4351 = ~new_G7417 | ~new_G7424;
  assign new_G4354 = ~new_G7425 | ~new_G7432;
  assign new_G4561 = ~new_G7518 | ~new_G7521;
  assign new_G4562 = ~new_G7515 | ~new_G7522;
  assign new_G4570 = ~new_G7526 | ~new_G7529;
  assign new_G4571 = ~new_G7523 | ~new_G7530;
  assign new_G4575 = ~new_G7554 | ~new_G7557;
  assign new_G4584 = ~new_G7562 | ~new_G7565;
  assign new_G4585 = ~new_G7559 | ~new_G7566;
  assign new_G4593 = ~new_G7570 | ~new_G7573;
  assign new_G4594 = ~new_G7567 | ~new_G7574;
  assign new_G4938 = ~new_G4929 | ~new_G4936;
  assign new_G4979 = ~new_G4970 | ~new_G4977;
  assign new_G6753 = ~new_G6748 | ~new_G6751;
  assign new_G6754 = ~new_G6745 | ~new_G6752;
  assign new_G6763 = ~new_G6758 | ~new_G6761;
  assign new_G6764 = ~new_G6755 | ~new_G6762;
  assign new_G6797 = ~new_G6792 | ~new_G6795;
  assign new_G6798 = ~new_G6789 | ~new_G6796;
  assign new_G6807 = ~new_G6802 | ~new_G6805;
  assign new_G6808 = ~new_G6799 | ~new_G6806;
  assign new_G7281 = ~new_G7276 | ~new_G7279;
  assign new_G7282 = ~new_G7273 | ~new_G7280;
  assign new_G7291 = ~new_G7286 | ~new_G7289;
  assign new_G7292 = ~new_G7283 | ~new_G7290;
  assign new_G7539 = ~new_G7534 | ~new_G7537;
  assign new_G7540 = ~new_G7531 | ~new_G7538;
  assign new_G7549 = ~new_G7544 | ~new_G7547;
  assign new_G7550 = ~new_G7541 | ~new_G7548;
  assign new_G7583 = ~new_G7578 | ~new_G7581;
  assign new_G7584 = ~new_G7575 | ~new_G7582;
  assign new_G7593 = ~new_G7588 | ~new_G7591;
  assign new_G7594 = ~new_G7585 | ~new_G7592;
  assign new_G1856 = ~new_G1850;
  assign new_G920 = new_G792 & new_G805 & new_G827 & new_G895 & new_G853;
  assign new_G925 = new_G792 & new_G821;
  assign new_G926 = new_G845 & new_G805 & new_G792;
  assign new_G927 = new_G805 & new_G868 & new_G827 & new_G792;
  assign new_G928 = new_G805 & new_G877 & new_G792 & new_G853 & new_G827;
  assign new_G937 = new_G805 & new_G845;
  assign new_G938 = new_G805 & new_G827 & new_G868;
  assign new_G939 = new_G805 & new_G877 & new_G853 & new_G827;
  assign new_G940 = new_G853 & new_G805 & new_G895 & new_G827;
  assign new_G941 = new_G805 & new_G845;
  assign new_G942 = new_G805 & new_G827 & new_G868;
  assign new_G943 = new_G805 & new_G877 & new_G853 & new_G827;
  assign new_G944 = new_G827 & new_G868;
  assign new_G945 = new_G877 & new_G853 & new_G827;
  assign new_G946 = new_G853 & new_G895 & new_G827;
  assign new_G947 = new_G827 & new_G868;
  assign new_G948 = new_G877 & new_G853 & new_G827;
  assign new_G949 = new_G853 & new_G877;
  assign new_G956 = new_G895 & new_G853;
  assign new_G1122 = new_G1074 & new_G1026 & new_G1055 & new_G1038 & new_G1093;
  assign new_G1125 = new_G1026 & new_G1050;
  assign new_G1126 = new_G1068 & new_G1038 & new_G1026;
  assign new_G1127 = new_G1038 & new_G1086 & new_G1055 & new_G1026;
  assign new_G1128 = new_G1038 & new_G1102 & new_G1026 & new_G1074 & new_G1055;
  assign new_G1132 = new_G1038 & new_G1068;
  assign new_G1133 = new_G1038 & new_G1055 & new_G1086;
  assign new_G1134 = new_G1038 & new_G1102 & new_G1074 & new_G1055;
  assign new_G1137 = new_G1086 & new_G1055;
  assign new_G1138 = new_G1102 & new_G1074 & new_G1055;
  assign new_G1141 = new_G1074 & new_G1102;
  assign new_G1221 = ~new_G1217;
  assign new_G1230 = ~new_G1226;
  assign new_G1244 = ~new_G1240;
  assign new_G1253 = ~new_G1249;
  assign new_G1267 = ~new_G1263;
  assign new_G1276 = ~new_G1272;
  assign new_G1284 = new_G1235;
  assign new_G1288 = new_G1235;
  assign new_G1292 = new_G1258;
  assign new_G1296 = new_G1258;
  assign new_G1300 = new_G1281;
  assign new_G1304 = new_G1281;
  assign new_G1702 = new_G1546 & new_G1556 & new_G1687 & new_G1573;
  assign new_G1705 = new_G1546 & new_G1567;
  assign new_G1706 = new_G1584 & new_G1556 & new_G1546;
  assign new_G1707 = new_G1556 & new_G1590 & new_G1573 & new_G1546;
  assign new_G1709 = new_G1556 & new_G1584;
  assign new_G1710 = new_G1556 & new_G1573 & new_G1590;
  assign new_G1711 = new_G1556 & new_G1687 & new_G1573;
  assign new_G1712 = new_G1556 & new_G1584;
  assign new_G1713 = new_G1556 & new_G1573 & new_G1590;
  assign new_G1714 = new_G1573 & new_G1590;
  assign new_G1718 = new_G1598 & new_G1609 & new_G1630 & new_G1695 & new_G1655;
  assign new_G1722 = new_G1598 & new_G1624;
  assign new_G1723 = new_G1647 & new_G1609 & new_G1598;
  assign new_G1724 = new_G1609 & new_G1669 & new_G1630 & new_G1598;
  assign new_G1725 = new_G1609 & new_G1677 & new_G1598 & new_G1655 & new_G1630;
  assign new_G1733 = new_G1609 & new_G1647;
  assign new_G1734 = new_G1609 & new_G1630 & new_G1669;
  assign new_G1735 = new_G1609 & new_G1677 & new_G1655 & new_G1630;
  assign new_G1736 = new_G1655 & new_G1609 & new_G1695 & new_G1630;
  assign new_G1737 = new_G1609 & new_G1647;
  assign new_G1738 = new_G1609 & new_G1630 & new_G1669;
  assign new_G1739 = new_G1609 & new_G1677 & new_G1655 & new_G1630;
  assign new_G1740 = new_G1630 & new_G1669;
  assign new_G1741 = new_G1677 & new_G1655 & new_G1630;
  assign new_G1742 = new_G1655 & new_G1695 & new_G1630;
  assign new_G1743 = new_G1630 & new_G1669;
  assign new_G1744 = new_G1677 & new_G1655 & new_G1630;
  assign new_G1745 = new_G1655 & new_G1677;
  assign new_G1749 = new_G1687 & new_G1573;
  assign new_G1750 = new_G1695 & new_G1655;
  assign new_G1935 = new_G1795 & new_G1822 & new_G1805 & new_G1850;
  assign new_G1938 = new_G1795 & new_G1816;
  assign new_G1939 = new_G1834 & new_G1805 & new_G1795;
  assign new_G1940 = new_G1805 & new_G1841 & new_G1822 & new_G1795;
  assign new_G1942 = new_G1805 & new_G1834;
  assign new_G1943 = new_G1805 & new_G1822 & new_G1841;
  assign new_G1944 = new_G1805 & new_G1850 & new_G1822;
  assign new_G1945 = new_G1805 & new_G1834;
  assign new_G1946 = new_G1805 & new_G1841 & new_G1822;
  assign new_G1947 = new_G1822 & new_G1841;
  assign new_G1948 = new_G1850 & new_G1822;
  assign new_G1949 = new_G1822 & new_G1841;
  assign new_G1950 = new_G1903 & new_G1859 & new_G1885 & new_G1869 & new_G1921;
  assign new_G1953 = new_G1859 & new_G1880;
  assign new_G1954 = new_G1897 & new_G1869 & new_G1859;
  assign new_G1955 = new_G1869 & new_G1914 & new_G1885 & new_G1859;
  assign new_G1956 = new_G1869 & new_G1929 & new_G1859 & new_G1903 & new_G1885;
  assign new_G1960 = new_G1869 & new_G1897;
  assign new_G1961 = new_G1869 & new_G1885 & new_G1914;
  assign new_G1962 = new_G1869 & new_G1929 & new_G1903 & new_G1885;
  assign new_G1965 = new_G1914 & new_G1885;
  assign new_G1966 = new_G1929 & new_G1903 & new_G1885;
  assign new_G1969 = new_G1903 & new_G1929;
  assign new_G2343 = ~new_G2341 | ~new_G2342;
  assign new_G2354 = ~new_G2352 | ~new_G2353;
  assign new_G2372 = ~new_G2370 | ~new_G2371;
  assign new_G2400 = ~new_G2398 | ~new_G2399;
  assign new_G2409 = ~new_G2407 | ~new_G2408;
  assign new_G2420 = ~new_G2418 | ~new_G2419;
  assign new_G2436 = ~new_G2434 | ~new_G2435;
  assign new_G2454 = ~new_G2452 | ~new_G2453;
  assign new_G2470 = ~new_G5932 | ~new_G5935;
  assign new_G5936 = ~new_G5932;
  assign new_G5983 = ~new_G5977;
  assign new_G2589 = ~new_G2587 | ~new_G2588;
  assign new_G2600 = ~new_G2598 | ~new_G2599;
  assign new_G2618 = ~new_G2616 | ~new_G2617;
  assign new_G2643 = ~new_G2641 | ~new_G2642;
  assign new_G2655 = ~new_G2653 | ~new_G2654;
  assign new_G2676 = ~new_G2674 | ~new_G2675;
  assign new_G2701 = ~new_G2699 | ~new_G2700;
  assign new_G2734 = ~new_G2732 | ~new_G2733;
  assign new_G2740 = ~new_G6052 | ~new_G6055;
  assign new_G6056 = ~new_G6052;
  assign new_G3022 = new_G2956 & new_G2965 & new_G3018 & new_G2973;
  assign new_G3025 = new_G2956 & new_G2970;
  assign new_G3026 = new_G2977 & new_G2965 & new_G2956;
  assign new_G3027 = new_G2965 & new_G2979 & new_G2973 & new_G2956;
  assign new_G3029 = new_G2982 & new_G2992 & new_G3001 & new_G3021 & new_G3009;
  assign new_G3030 = new_G2982 & new_G2998;
  assign new_G3031 = new_G3006 & new_G2992 & new_G2982;
  assign new_G3032 = new_G2992 & new_G3013 & new_G3001 & new_G2982;
  assign new_G3033 = new_G2992 & new_G3015 & new_G2982 & new_G3009 & new_G3001;
  assign new_G3052 = ~new_G3050 | ~new_G3051;
  assign new_G3062 = ~new_G3060 | ~new_G3061;
  assign new_G3071 = ~new_G3069 | ~new_G3070;
  assign new_G3082 = ~new_G3080 | ~new_G3081;
  assign new_G3093 = ~new_G3091 | ~new_G3092;
  assign new_G3102 = ~new_G3100 | ~new_G3101;
  assign new_G3110 = ~new_G3108 | ~new_G3109;
  assign new_G3119 = ~new_G3117 | ~new_G3118;
  assign new_G3122 = ~new_G3120 | ~new_G3121;
  assign new_G3228 = new_G3176 & new_G3186 & new_G3195 & new_G3215 & new_G3203;
  assign new_G3231 = new_G3176 & new_G3192;
  assign new_G3232 = new_G3200 & new_G3186 & new_G3176;
  assign new_G3233 = new_G3186 & new_G3207 & new_G3195 & new_G3176;
  assign new_G3234 = new_G3186 & new_G3209 & new_G3176 & new_G3203 & new_G3195;
  assign new_G3283 = ~new_G3281 | ~new_G3282;
  assign new_G3295 = ~new_G3293 | ~new_G3294;
  assign new_G3314 = ~new_G3312 | ~new_G3313;
  assign new_G3344 = ~new_G3342 | ~new_G3343;
  assign new_G3353 = ~new_G3351 | ~new_G3352;
  assign new_G3365 = ~new_G3363 | ~new_G3364;
  assign new_G3381 = ~new_G3379 | ~new_G3380;
  assign new_G3399 = ~new_G3397 | ~new_G3398;
  assign new_G3417 = ~new_G3415 | ~new_G3416;
  assign new_G6685 = ~new_G6679;
  assign new_G3508 = ~new_G3504;
  assign new_G3517 = ~new_G3513;
  assign new_G3527 = ~new_G3525 | ~new_G3526;
  assign new_G3536 = ~new_G3534 | ~new_G3535;
  assign new_G3545 = ~new_G3543 | ~new_G3544;
  assign new_G3550 = ~new_G3548 | ~new_G3549;
  assign new_G3559 = ~new_G3557 | ~new_G3558;
  assign new_G3568 = ~new_G3566 | ~new_G3567;
  assign new_G3571 = new_G3522;
  assign new_G3575 = new_G3522;
  assign new_G3845 = ~new_G3843 | ~new_G3844;
  assign new_G3856 = ~new_G3854 | ~new_G3855;
  assign new_G3874 = ~new_G3872 | ~new_G3873;
  assign new_G3899 = ~new_G3897 | ~new_G3898;
  assign new_G3911 = ~new_G3909 | ~new_G3910;
  assign new_G3932 = ~new_G3930 | ~new_G3931;
  assign new_G3957 = ~new_G3955 | ~new_G3956;
  assign new_G3989 = ~new_G3987 | ~new_G3988;
  assign new_G3997 = ~new_G3995 | ~new_G3996;
  assign new_G4180 = ~new_G4178 | ~new_G4179;
  assign new_G4189 = ~new_G4187 | ~new_G4188;
  assign new_G4198 = ~new_G4196 | ~new_G4197;
  assign new_G4207 = ~new_G4203;
  assign new_G4216 = ~new_G4212;
  assign new_G4221 = ~new_G4219 | ~new_G4220;
  assign new_G4230 = ~new_G4226;
  assign new_G4239 = ~new_G4235;
  assign new_G4263 = new_G4244;
  assign new_G4267 = new_G4244;
  assign new_G4291 = ~new_G4289 | ~new_G4290;
  assign new_G4300 = ~new_G4298 | ~new_G4299;
  assign new_G4308 = ~new_G4306 | ~new_G4307;
  assign new_G4317 = ~new_G4315 | ~new_G4316;
  assign new_G4327 = ~new_G4325 | ~new_G4326;
  assign new_G4336 = ~new_G4334 | ~new_G4335;
  assign new_G4344 = ~new_G4342 | ~new_G4343;
  assign new_G4352 = ~new_G4350 | ~new_G4351;
  assign new_G4355 = ~new_G4353 | ~new_G4354;
  assign new_G4535 = ~new_G4531;
  assign new_G4544 = ~new_G4540;
  assign new_G4558 = ~new_G4554;
  assign new_G4563 = ~new_G4561 | ~new_G4562;
  assign new_G4572 = ~new_G4570 | ~new_G4571;
  assign new_G4577 = ~new_G4575 | ~new_G4576;
  assign new_G4586 = ~new_G4584 | ~new_G4585;
  assign new_G4595 = ~new_G4593 | ~new_G4594;
  assign new_G4598 = new_G4549;
  assign new_G4602 = new_G4549;
  assign new_G4716 = new_G1921;
  assign new_G4724 = new_G1859;
  assign new_G4732 = new_G1869;
  assign new_G4740 = new_G1885;
  assign new_G4748 = new_G1903;
  assign new_G4756 = new_G1093;
  assign new_G4764 = new_G1026;
  assign new_G4772 = new_G1038;
  assign new_G4780 = new_G1055;
  assign new_G4788 = new_G1074;
  assign new_G4939 = ~new_G4937 | ~new_G4938;
  assign new_G4980 = ~new_G4978 | ~new_G4979;
  assign new_G5044 = new_G895;
  assign new_G5054 = new_G853;
  assign new_G5064 = new_G792;
  assign new_G5074 = new_G827;
  assign new_G5084 = new_G805;
  assign new_G5094 = new_G805;
  assign new_G5132 = new_G895;
  assign new_G5142 = new_G853;
  assign new_G5152 = new_G792;
  assign new_G5162 = new_G827;
  assign new_G5365 = ~new_G5359;
  assign new_G5366 = ~new_G5362;
  assign new_G5488 = new_G1687;
  assign new_G5498 = new_G1573;
  assign new_G5508 = new_G1546;
  assign new_G5518 = new_G1556;
  assign new_G5546 = new_G1687;
  assign new_G5556 = new_G1573;
  assign new_G5566 = new_G1546;
  assign new_G5576 = new_G1556;
  assign new_G5614 = new_G1695;
  assign new_G5624 = new_G1655;
  assign new_G5634 = new_G1598;
  assign new_G5644 = new_G1630;
  assign new_G5654 = new_G1609;
  assign new_G5664 = new_G1609;
  assign new_G5702 = new_G1695;
  assign new_G5712 = new_G1655;
  assign new_G5722 = new_G1598;
  assign new_G5732 = new_G1630;
  assign new_G5820 = new_G1795;
  assign new_G5828 = new_G1795;
  assign new_G5836 = new_G1805;
  assign new_G5844 = new_G1805;
  assign new_G5852 = new_G1822;
  assign new_G5860 = new_G1822;
  assign new_G6121 = ~new_G6115;
  assign new_G6179 = ~new_G6173;
  assign new_G6261 = new_G2724;
  assign new_G7359 = ~new_G7353;
  assign new_G7360 = ~new_G7356;
  assign new_G7343 = ~new_G7337;
  assign new_G7344 = ~new_G7340;
  assign new_G6809 = ~new_G6763 | ~new_G6764;
  assign new_G6812 = ~new_G6753 | ~new_G6754;
  assign new_G6819 = ~new_G6807 | ~new_G6808;
  assign new_G6822 = ~new_G6797 | ~new_G6798;
  assign new_G6989 = ~new_G6983;
  assign new_G7135 = ~new_G7129;
  assign new_G7345 = ~new_G7291 | ~new_G7292;
  assign new_G7348 = ~new_G7281 | ~new_G7282;
  assign new_G7601 = ~new_G7595;
  assign new_G7602 = ~new_G7598;
  assign new_G7603 = ~new_G7549 | ~new_G7550;
  assign new_G7606 = ~new_G7539 | ~new_G7540;
  assign new_G7611 = ~new_G7593 | ~new_G7594;
  assign new_G7614 = ~new_G7583 | ~new_G7584;
  assign new_G929 = new_G928 | new_G927 | new_G926 | new_G802 | new_G925;
  assign new_G950 = new_G868 | new_G949;
  assign new_G1129 = new_G1128 | new_G1127 | new_G1126 | new_G1035 | new_G1125;
  assign new_G1708 = new_G1707 | new_G1706 | new_G1553 | new_G1705;
  assign new_G1715 = new_G1584 | new_G1714;
  assign new_G1726 = new_G1725 | new_G1724 | new_G1723 | new_G1606 | new_G1722;
  assign new_G1746 = new_G1669 | new_G1745;
  assign new_G1941 = new_G1940 | new_G1939 | new_G1802 | new_G1938;
  assign new_G1957 = new_G1956 | new_G1955 | new_G1954 | new_G1866 | new_G1953;
  assign new_G2471 = ~new_G5929 | ~new_G5936;
  assign new_G2741 = ~new_G6049 | ~new_G6056;
  assign new_G3028 = new_G3027 | new_G3026 | new_G2962 | new_G3025;
  assign new_G3034 = new_G3033 | new_G3032 | new_G3031 | new_G2989 | new_G3030;
  assign new_G3235 = new_G3234 | new_G3233 | new_G3232 | new_G3183 | new_G3231;
  assign new_G5014 = new_G946 | new_G945 | new_G845 | new_G944;
  assign new_G5034 = new_G940 | new_G939 | new_G938 | new_G821 | new_G937;
  assign new_G5102 = ~new_G948 & ~new_G845 & ~new_G947;
  assign new_G5122 = ~new_G943 & ~new_G942 & ~new_G821 & ~new_G941;
  assign new_G5367 = ~new_G5362 | ~new_G5365;
  assign new_G5368 = ~new_G5359 | ~new_G5366;
  assign new_G5478 = new_G1711 | new_G1710 | new_G1567 | new_G1709;
  assign new_G5536 = ~new_G1713 & ~new_G1567 & ~new_G1712;
  assign new_G5584 = new_G1742 | new_G1741 | new_G1647 | new_G1740;
  assign new_G5604 = new_G1736 | new_G1735 | new_G1734 | new_G1624 | new_G1733;
  assign new_G5672 = ~new_G1744 & ~new_G1647 & ~new_G1743;
  assign new_G5692 = ~new_G1739 & ~new_G1738 & ~new_G1624 & ~new_G1737;
  assign new_G5817 = new_G1944 | new_G1943 | new_G1816 | new_G1942;
  assign new_G5825 = ~new_G1946 & ~new_G1816 & ~new_G1945;
  assign new_G5833 = new_G1948 | new_G1834 | new_G1947;
  assign new_G5841 = ~new_G1834 & ~new_G1949;
  assign new_G6340 = ~new_G7356 | ~new_G7359;
  assign new_G6341 = ~new_G7353 | ~new_G7360;
  assign new_G6350 = ~new_G7340 | ~new_G7343;
  assign new_G6351 = ~new_G7337 | ~new_G7344;
  assign new_G7436 = ~new_G7598 | ~new_G7601;
  assign new_G7437 = ~new_G7595 | ~new_G7602;
  assign new_G4720 = ~new_G4716;
  assign new_G4728 = ~new_G4724;
  assign new_G4736 = ~new_G4732;
  assign new_G4744 = ~new_G4740;
  assign new_G4752 = ~new_G4748;
  assign new_G4760 = ~new_G4756;
  assign new_G4768 = ~new_G4764;
  assign new_G4776 = ~new_G4772;
  assign new_G4784 = ~new_G4780;
  assign new_G4792 = ~new_G4788;
  assign new_G3350 = ~new_G3344;
  assign new_G2406 = ~new_G2400;
  assign new_G924 = ~new_G920;
  assign new_G5088 = ~new_G5084;
  assign new_G5098 = ~new_G5094;
  assign new_G997 = new_G902 & new_G920;
  assign new_G1146 = new_G1108 & new_G1122;
  assign new_G1287 = ~new_G1284;
  assign new_G1291 = ~new_G1288;
  assign new_G1295 = ~new_G1292;
  assign new_G1299 = ~new_G1296;
  assign new_G1303 = ~new_G1300;
  assign new_G1307 = ~new_G1304;
  assign new_G1309 = new_G1284 & new_G1226 & new_G1217;
  assign new_G1312 = new_G1288 & new_G1230 & new_G1221;
  assign new_G1315 = new_G1292 & new_G1249 & new_G1240;
  assign new_G1318 = new_G1296 & new_G1253 & new_G1244;
  assign new_G1321 = new_G1300 & new_G1272 & new_G1263;
  assign new_G1324 = new_G1304 & new_G1276 & new_G1267;
  assign new_G1721 = ~new_G1718;
  assign new_G5522 = ~new_G5518;
  assign new_G5580 = ~new_G5576;
  assign new_G5658 = ~new_G5654;
  assign new_G5668 = ~new_G5664;
  assign new_G1788 = new_G1702 & new_G1718;
  assign new_G1974 = new_G1935 & new_G1950;
  assign new_G5824 = ~new_G5820;
  assign new_G5832 = ~new_G5828;
  assign new_G5840 = ~new_G5836;
  assign new_G5848 = ~new_G5844;
  assign new_G1999 = ~new_G5852 | ~new_G5855;
  assign new_G5856 = ~new_G5852;
  assign new_G2003 = ~new_G5860 | ~new_G5863;
  assign new_G5864 = ~new_G5860;
  assign new_G2472 = ~new_G2470 | ~new_G2471;
  assign new_G2487 = new_G2343 & new_G2372 & new_G2354 & new_G2400;
  assign new_G2492 = new_G2343 & new_G2366;
  assign new_G2493 = new_G2384 & new_G2354 & new_G2343;
  assign new_G2494 = new_G2354 & new_G2391 & new_G2372 & new_G2343;
  assign new_G2500 = new_G2354 & new_G2384;
  assign new_G2501 = new_G2354 & new_G2372 & new_G2391;
  assign new_G2502 = new_G2354 & new_G2400 & new_G2372;
  assign new_G2503 = new_G2354 & new_G2384;
  assign new_G2504 = new_G2354 & new_G2391 & new_G2372;
  assign new_G2505 = new_G2372 & new_G2391;
  assign new_G2506 = new_G2400 & new_G2372;
  assign new_G2507 = new_G2372 & new_G2391;
  assign new_G2511 = new_G2409 & new_G2431;
  assign new_G2512 = new_G2448 & new_G2420 & new_G2409;
  assign new_G2513 = new_G2420 & new_G2465 & new_G2436 & new_G2409;
  assign new_G2514 = new_G2420 & new_G2481 & new_G2409 & new_G2454 & new_G2436;
  assign new_G2518 = new_G2420 & new_G2448;
  assign new_G2519 = new_G2420 & new_G2436 & new_G2465;
  assign new_G2520 = new_G2420 & new_G2481 & new_G2454 & new_G2436;
  assign new_G2523 = new_G2465 & new_G2436;
  assign new_G2524 = new_G2481 & new_G2454 & new_G2436;
  assign new_G2527 = new_G2454 & new_G2481;
  assign new_G2742 = ~new_G2740 | ~new_G2741;
  assign new_G2749 = new_G2589 & new_G2600 & new_G2734 & new_G2618;
  assign new_G2754 = new_G2589 & new_G2612;
  assign new_G2755 = new_G2629 & new_G2600 & new_G2589;
  assign new_G2756 = new_G2600 & new_G2635 & new_G2618 & new_G2589;
  assign new_G2762 = new_G2600 & new_G2629;
  assign new_G2763 = new_G2600 & new_G2618 & new_G2635;
  assign new_G2764 = new_G2600 & new_G2734 & new_G2618;
  assign new_G2765 = new_G2600 & new_G2629;
  assign new_G2766 = new_G2600 & new_G2618 & new_G2635;
  assign new_G2767 = new_G2618 & new_G2635;
  assign new_G2776 = new_G2643 & new_G2670;
  assign new_G2777 = new_G2693 & new_G2655 & new_G2643;
  assign new_G2778 = new_G2655 & new_G2715 & new_G2676 & new_G2643;
  assign new_G2779 = new_G2655 & new_G2724 & new_G2643 & new_G2701 & new_G2676;
  assign new_G2788 = new_G2655 & new_G2693;
  assign new_G2789 = new_G2655 & new_G2676 & new_G2715;
  assign new_G2790 = new_G2655 & new_G2724 & new_G2701 & new_G2676;
  assign new_G2792 = new_G2655 & new_G2693;
  assign new_G2793 = new_G2655 & new_G2676 & new_G2715;
  assign new_G2794 = new_G2655 & new_G2724 & new_G2701 & new_G2676;
  assign new_G2795 = new_G2676 & new_G2715;
  assign new_G2796 = new_G2724 & new_G2701 & new_G2676;
  assign new_G2798 = new_G2676 & new_G2715;
  assign new_G2799 = new_G2724 & new_G2701 & new_G2676;
  assign new_G2800 = new_G2701 & new_G2724;
  assign new_G2804 = new_G2734 & new_G2618;
  assign new_G3035 = new_G3022 & new_G3029;
  assign new_G3045 = new_G3022 & new_G3034;
  assign new_G3123 = new_G3052 & new_G3062 & new_G3119 & new_G3071;
  assign new_G3128 = new_G3052 & new_G3068;
  assign new_G3129 = new_G3076 & new_G3062 & new_G3052;
  assign new_G3130 = new_G3062 & new_G3079 & new_G3071 & new_G3052;
  assign new_G3136 = new_G3082 & new_G3093 & new_G3102 & new_G3122 & new_G3110;
  assign new_G3139 = new_G3082 & new_G3099;
  assign new_G3140 = new_G3107 & new_G3093 & new_G3082;
  assign new_G3141 = new_G3093 & new_G3114 & new_G3102 & new_G3082;
  assign new_G3142 = new_G3093 & new_G3116 & new_G3082 & new_G3110 & new_G3102;
  assign new_G3249 = new_G3216 & new_G3228;
  assign new_G3431 = new_G3283 & new_G3314 & new_G3295 & new_G3344;
  assign new_G3434 = new_G3283 & new_G3308;
  assign new_G3435 = new_G3327 & new_G3295 & new_G3283;
  assign new_G3436 = new_G3295 & new_G3335 & new_G3314 & new_G3283;
  assign new_G3438 = new_G3295 & new_G3327;
  assign new_G3439 = new_G3295 & new_G3314 & new_G3335;
  assign new_G3440 = new_G3295 & new_G3344 & new_G3314;
  assign new_G3441 = new_G3295 & new_G3327;
  assign new_G3442 = new_G3295 & new_G3335 & new_G3314;
  assign new_G3443 = new_G3314 & new_G3335;
  assign new_G3444 = new_G3344 & new_G3314;
  assign new_G3445 = new_G3314 & new_G3335;
  assign new_G3446 = new_G3399 & new_G3353 & new_G3381 & new_G3365 & new_G3417;
  assign new_G3449 = new_G3353 & new_G3376;
  assign new_G3450 = new_G3393 & new_G3365 & new_G3353;
  assign new_G3451 = new_G3365 & new_G3410 & new_G3381 & new_G3353;
  assign new_G3452 = new_G3365 & new_G3425 & new_G3353 & new_G3399 & new_G3381;
  assign new_G3456 = new_G3365 & new_G3393;
  assign new_G3457 = new_G3365 & new_G3381 & new_G3410;
  assign new_G3458 = new_G3365 & new_G3425 & new_G3399 & new_G3381;
  assign new_G3460 = new_G3410 & new_G3381;
  assign new_G3461 = new_G3425 & new_G3399 & new_G3381;
  assign new_G3463 = new_G3399 & new_G3425;
  assign new_G3531 = ~new_G3527;
  assign new_G3540 = ~new_G3536;
  assign new_G3554 = ~new_G3550;
  assign new_G3563 = ~new_G3559;
  assign new_G3574 = ~new_G3571;
  assign new_G3578 = ~new_G3575;
  assign new_G3579 = new_G3545;
  assign new_G3583 = new_G3545;
  assign new_G3587 = new_G3568;
  assign new_G3591 = new_G3568;
  assign new_G3596 = new_G3571 & new_G3513 & new_G3504;
  assign new_G3599 = new_G3575 & new_G3517 & new_G3508;
  assign new_G4004 = new_G3845 & new_G3856 & new_G3989 & new_G3874;
  assign new_G4007 = new_G3845 & new_G3868;
  assign new_G4008 = new_G3885 & new_G3856 & new_G3845;
  assign new_G4009 = new_G3856 & new_G3891 & new_G3874 & new_G3845;
  assign new_G4011 = new_G3856 & new_G3885;
  assign new_G4012 = new_G3856 & new_G3874 & new_G3891;
  assign new_G4013 = new_G3856 & new_G3989 & new_G3874;
  assign new_G4014 = new_G3856 & new_G3885;
  assign new_G4015 = new_G3856 & new_G3874 & new_G3891;
  assign new_G4016 = new_G3874 & new_G3891;
  assign new_G4020 = new_G3899 & new_G3911 & new_G3932 & new_G3997 & new_G3957;
  assign new_G4024 = new_G3899 & new_G3926;
  assign new_G4025 = new_G3949 & new_G3911 & new_G3899;
  assign new_G4026 = new_G3911 & new_G3971 & new_G3932 & new_G3899;
  assign new_G4027 = new_G3911 & new_G3979 & new_G3899 & new_G3957 & new_G3932;
  assign new_G4035 = new_G3911 & new_G3949;
  assign new_G4036 = new_G3911 & new_G3932 & new_G3971;
  assign new_G4037 = new_G3911 & new_G3979 & new_G3957 & new_G3932;
  assign new_G4038 = new_G3957 & new_G3911 & new_G3997 & new_G3932;
  assign new_G4039 = new_G3911 & new_G3949;
  assign new_G4040 = new_G3911 & new_G3932 & new_G3971;
  assign new_G4041 = new_G3911 & new_G3979 & new_G3957 & new_G3932;
  assign new_G4042 = new_G3932 & new_G3971;
  assign new_G4043 = new_G3979 & new_G3957 & new_G3932;
  assign new_G4044 = new_G3957 & new_G3997 & new_G3932;
  assign new_G4045 = new_G3932 & new_G3971;
  assign new_G4046 = new_G3979 & new_G3957 & new_G3932;
  assign new_G4047 = new_G3957 & new_G3979;
  assign new_G4051 = new_G3989 & new_G3874;
  assign new_G4052 = new_G3997 & new_G3957;
  assign new_G4184 = ~new_G4180;
  assign new_G4193 = ~new_G4189;
  assign new_G4247 = new_G4198;
  assign new_G4251 = new_G4198;
  assign new_G4255 = new_G4221;
  assign new_G4259 = new_G4221;
  assign new_G4266 = ~new_G4263;
  assign new_G4270 = ~new_G4267;
  assign new_G4284 = new_G4263 & new_G4235 & new_G4226;
  assign new_G4287 = new_G4267 & new_G4239 & new_G4230;
  assign new_G4356 = new_G4291 & new_G4300 & new_G4352 & new_G4308;
  assign new_G4361 = new_G4291 & new_G4305;
  assign new_G4362 = new_G4312 & new_G4300 & new_G4291;
  assign new_G4363 = new_G4300 & new_G4314 & new_G4308 & new_G4291;
  assign new_G4369 = new_G4317 & new_G4327 & new_G4336 & new_G4355 & new_G4344;
  assign new_G4372 = new_G4317 & new_G4333;
  assign new_G4373 = new_G4341 & new_G4327 & new_G4317;
  assign new_G4374 = new_G4327 & new_G4348 & new_G4336 & new_G4317;
  assign new_G4375 = new_G4327 & new_G4349 & new_G4317 & new_G4344 & new_G4336;
  assign new_G4567 = ~new_G4563;
  assign new_G4581 = ~new_G4577;
  assign new_G4590 = ~new_G4586;
  assign new_G4601 = ~new_G4598;
  assign new_G4605 = ~new_G4602;
  assign new_G4606 = new_G4572;
  assign new_G4610 = new_G4572;
  assign new_G4614 = new_G4595;
  assign new_G4618 = new_G4595;
  assign new_G4623 = new_G4598 & new_G4540 & new_G4531;
  assign new_G4626 = new_G4602 & new_G4544 & new_G4535;
  assign new_G4796 = new_G3417;
  assign new_G4804 = new_G3353;
  assign new_G4812 = new_G3365;
  assign new_G4820 = new_G3381;
  assign new_G4828 = new_G3399;
  assign new_G4844 = new_G2409;
  assign new_G4852 = new_G2420;
  assign new_G4860 = new_G2436;
  assign new_G4868 = new_G2454;
  assign new_G4945 = ~new_G4939;
  assign new_G4948 = ~new_G4939 | ~new_G4946;
  assign new_G4986 = ~new_G4980;
  assign new_G4989 = ~new_G4980 | ~new_G4987;
  assign new_G5048 = ~new_G5044;
  assign new_G5058 = ~new_G5054;
  assign new_G5068 = ~new_G5064;
  assign new_G5078 = ~new_G5074;
  assign new_G5166 = ~new_G5162;
  assign new_G5136 = ~new_G5132;
  assign new_G5146 = ~new_G5142;
  assign new_G5156 = ~new_G5152;
  assign new_G5388 = ~new_G5367 | ~new_G5368;
  assign new_G5492 = ~new_G5488;
  assign new_G5502 = ~new_G5498;
  assign new_G5512 = ~new_G5508;
  assign new_G5550 = ~new_G5546;
  assign new_G5560 = ~new_G5556;
  assign new_G5570 = ~new_G5566;
  assign new_G5618 = ~new_G5614;
  assign new_G5628 = ~new_G5624;
  assign new_G5638 = ~new_G5634;
  assign new_G5648 = ~new_G5644;
  assign new_G5736 = ~new_G5732;
  assign new_G5706 = ~new_G5702;
  assign new_G5716 = ~new_G5712;
  assign new_G5726 = ~new_G5722;
  assign new_G5940 = new_G2343;
  assign new_G5948 = new_G2343;
  assign new_G5956 = new_G2354;
  assign new_G5964 = new_G2354;
  assign new_G5972 = new_G2372;
  assign new_G5980 = new_G2372;
  assign new_G6080 = new_G2734;
  assign new_G6090 = new_G2618;
  assign new_G6100 = new_G2589;
  assign new_G6110 = new_G2600;
  assign new_G6138 = new_G2734;
  assign new_G6148 = new_G2618;
  assign new_G6158 = new_G2589;
  assign new_G6168 = new_G2600;
  assign new_G6216 = new_G2701;
  assign new_G6226 = new_G2643;
  assign new_G6236 = new_G2676;
  assign new_G6246 = new_G2655;
  assign new_G6256 = new_G2655;
  assign new_G6267 = ~new_G6261;
  assign new_G6304 = new_G2701;
  assign new_G6314 = new_G2643;
  assign new_G6324 = new_G2676;
  assign new_G6342 = ~new_G6340 | ~new_G6341;
  assign new_G6352 = ~new_G6350 | ~new_G6351;
  assign new_G7351 = ~new_G7345;
  assign new_G7352 = ~new_G7348;
  assign new_G6642 = new_G3283;
  assign new_G6650 = new_G3283;
  assign new_G6658 = new_G3295;
  assign new_G6666 = new_G3295;
  assign new_G6674 = new_G3314;
  assign new_G6682 = new_G3314;
  assign new_G6815 = ~new_G6809;
  assign new_G6816 = ~new_G6812;
  assign new_G6825 = ~new_G6819;
  assign new_G6826 = ~new_G6822;
  assign new_G6948 = new_G3989;
  assign new_G6958 = new_G3874;
  assign new_G6968 = new_G3845;
  assign new_G6978 = new_G3856;
  assign new_G7006 = new_G3989;
  assign new_G7016 = new_G3874;
  assign new_G7026 = new_G3845;
  assign new_G7036 = new_G3856;
  assign new_G7074 = new_G3997;
  assign new_G7084 = new_G3957;
  assign new_G7094 = new_G3899;
  assign new_G7104 = new_G3932;
  assign new_G7114 = new_G3911;
  assign new_G7124 = new_G3911;
  assign new_G7162 = new_G3997;
  assign new_G7172 = new_G3957;
  assign new_G7182 = new_G3899;
  assign new_G7192 = new_G3932;
  assign new_G7438 = ~new_G7436 | ~new_G7437;
  assign new_G7617 = ~new_G7611;
  assign new_G7618 = ~new_G7614;
  assign new_G7609 = ~new_G7603;
  assign new_G7610 = ~new_G7606;
  assign new_G1151 = new_G1129 & new_G1108;
  assign new_G1002 = new_G902 & new_G929;
  assign new_G933 = ~new_G929;
  assign new_G1308 = new_G1287 & new_G1221 & new_G1226;
  assign new_G1311 = new_G1291 & new_G1217 & new_G1230;
  assign new_G1314 = new_G1295 & new_G1244 & new_G1249;
  assign new_G1317 = new_G1299 & new_G1240 & new_G1253;
  assign new_G1320 = new_G1303 & new_G1267 & new_G1272;
  assign new_G1323 = new_G1307 & new_G1263 & new_G1276;
  assign new_G1730 = ~new_G1726;
  assign new_G1789 = new_G1702 & new_G1726;
  assign new_G1981 = new_G1957 & new_G1935;
  assign new_G5823 = ~new_G5817;
  assign new_G1986 = ~new_G5817 | ~new_G5824;
  assign new_G5831 = ~new_G5825;
  assign new_G1989 = ~new_G5825 | ~new_G5832;
  assign new_G5839 = ~new_G5833;
  assign new_G1993 = ~new_G5833 | ~new_G5840;
  assign new_G5847 = ~new_G5841;
  assign new_G1996 = ~new_G5841 | ~new_G5848;
  assign new_G2000 = ~new_G5849 | ~new_G5856;
  assign new_G2004 = ~new_G5857 | ~new_G5864;
  assign new_G2495 = new_G2494 | new_G2493 | new_G2351 | new_G2492;
  assign new_G2515 = new_G2514 | new_G2513 | new_G2512 | new_G2417 | new_G2511;
  assign new_G2757 = new_G2756 | new_G2755 | new_G2597 | new_G2754;
  assign new_G2768 = new_G2629 | new_G2767;
  assign new_G2780 = new_G2779 | new_G2778 | new_G2777 | new_G2652 | new_G2776;
  assign new_G2801 = new_G2715 | new_G2800;
  assign new_G3046 = new_G3028 | new_G3045;
  assign new_G3131 = new_G3130 | new_G3129 | new_G3059 | new_G3128;
  assign new_G3143 = new_G3142 | new_G3141 | new_G3140 | new_G3090 | new_G3139;
  assign new_G3238 = ~new_G3235;
  assign new_G3258 = new_G3216 & new_G3235;
  assign new_G3437 = new_G3436 | new_G3435 | new_G3292 | new_G3434;
  assign new_G3453 = new_G3452 | new_G3451 | new_G3450 | new_G3362 | new_G3449;
  assign new_G3595 = new_G3574 & new_G3508 & new_G3513;
  assign new_G3598 = new_G3578 & new_G3504 & new_G3517;
  assign new_G4010 = new_G4009 | new_G4008 | new_G3853 | new_G4007;
  assign new_G4017 = new_G3885 | new_G4016;
  assign new_G4028 = new_G4027 | new_G4026 | new_G4025 | new_G3908 | new_G4024;
  assign new_G4048 = new_G3971 | new_G4047;
  assign new_G4283 = new_G4266 & new_G4230 & new_G4235;
  assign new_G4286 = new_G4270 & new_G4226 & new_G4239;
  assign new_G4364 = new_G4363 | new_G4362 | new_G4297 | new_G4361;
  assign new_G4376 = new_G4375 | new_G4374 | new_G4373 | new_G4324 | new_G4372;
  assign new_G4622 = new_G4601 & new_G4535 & new_G4540;
  assign new_G4625 = new_G4605 & new_G4531 & new_G4544;
  assign new_G4947 = ~new_G4942 | ~new_G4945;
  assign new_G4988 = ~new_G4983 | ~new_G4986;
  assign new_G5018 = ~new_G5014;
  assign new_G5019 = ~new_G5014 | ~new_G5017;
  assign new_G5024 = new_G950 | new_G956;
  assign new_G5038 = ~new_G5034;
  assign new_G5106 = ~new_G5102;
  assign new_G5107 = ~new_G5102 | ~new_G5105;
  assign new_G5112 = ~new_G950;
  assign new_G5126 = ~new_G5122;
  assign new_G5468 = new_G1715 | new_G1749;
  assign new_G5482 = ~new_G5478;
  assign new_G5526 = ~new_G1715;
  assign new_G5540 = ~new_G5536;
  assign new_G5588 = ~new_G5584;
  assign new_G5589 = ~new_G5584 | ~new_G5587;
  assign new_G5594 = new_G1746 | new_G1750;
  assign new_G5608 = ~new_G5604;
  assign new_G5676 = ~new_G5672;
  assign new_G5677 = ~new_G5672 | ~new_G5675;
  assign new_G5682 = ~new_G1746;
  assign new_G5696 = ~new_G5692;
  assign new_G5937 = new_G2502 | new_G2501 | new_G2366 | new_G2500;
  assign new_G5945 = ~new_G2504 & ~new_G2366 & ~new_G2503;
  assign new_G5953 = new_G2506 | new_G2384 | new_G2505;
  assign new_G5961 = ~new_G2384 & ~new_G2507;
  assign new_G6070 = new_G2764 | new_G2763 | new_G2612 | new_G2762;
  assign new_G6128 = ~new_G2766 & ~new_G2612 & ~new_G2765;
  assign new_G6264 = ~new_G2799 & ~new_G2693 & ~new_G2798;
  assign new_G6284 = ~new_G2794 & ~new_G2793 & ~new_G2670 & ~new_G2792;
  assign new_G6360 = ~new_G7348 | ~new_G7351;
  assign new_G6361 = ~new_G7345 | ~new_G7352;
  assign new_G6639 = new_G3440 | new_G3439 | new_G3308 | new_G3438;
  assign new_G6647 = ~new_G3442 & ~new_G3308 & ~new_G3441;
  assign new_G6655 = new_G3444 | new_G3327 | new_G3443;
  assign new_G6663 = ~new_G3327 & ~new_G3445;
  assign new_G6817 = ~new_G6812 | ~new_G6815;
  assign new_G6818 = ~new_G6809 | ~new_G6816;
  assign new_G6827 = ~new_G6822 | ~new_G6825;
  assign new_G6828 = ~new_G6819 | ~new_G6826;
  assign new_G6938 = new_G4013 | new_G4012 | new_G3868 | new_G4011;
  assign new_G6996 = ~new_G4015 & ~new_G3868 & ~new_G4014;
  assign new_G7044 = new_G4044 | new_G4043 | new_G3949 | new_G4042;
  assign new_G7064 = new_G4038 | new_G4037 | new_G4036 | new_G3926 | new_G4035;
  assign new_G7132 = ~new_G4046 & ~new_G3949 & ~new_G4045;
  assign new_G7152 = ~new_G4041 & ~new_G4040 & ~new_G3926 & ~new_G4039;
  assign new_G7446 = ~new_G7614 | ~new_G7617;
  assign new_G7447 = ~new_G7611 | ~new_G7618;
  assign new_G7456 = ~new_G7606 | ~new_G7609;
  assign new_G7457 = ~new_G7603 | ~new_G7610;
  assign new_G241 = new_G1117 | new_G1151;
  assign new_G265 = new_G908 | new_G1002;
  assign new_G2005 = ~new_G2003 | ~new_G2004;
  assign new_G4800 = ~new_G4796;
  assign new_G4808 = ~new_G4804;
  assign new_G4816 = ~new_G4812;
  assign new_G4824 = ~new_G4820;
  assign new_G4832 = ~new_G4828;
  assign new_G4848 = ~new_G4844;
  assign new_G4856 = ~new_G4852;
  assign new_G4864 = ~new_G4860;
  assign new_G4872 = ~new_G4868;
  assign new_G1310 = ~new_G1308 & ~new_G1309;
  assign new_G1313 = ~new_G1311 & ~new_G1312;
  assign new_G1316 = ~new_G1314 & ~new_G1315;
  assign new_G1319 = ~new_G1317 & ~new_G1318;
  assign new_G1322 = ~new_G1320 & ~new_G1321;
  assign new_G1325 = ~new_G1323 & ~new_G1324;
  assign new_G5392 = ~new_G5388;
  assign new_G1790 = new_G1708 | new_G1789;
  assign new_G1982 = new_G1941 | new_G1981;
  assign new_G1985 = ~new_G5820 | ~new_G5823;
  assign new_G1988 = ~new_G5828 | ~new_G5831;
  assign new_G1992 = ~new_G5836 | ~new_G5839;
  assign new_G1995 = ~new_G5844 | ~new_G5847;
  assign new_G2001 = ~new_G1999 | ~new_G2000;
  assign new_G2491 = ~new_G2487;
  assign new_G2508 = new_G2454 & new_G2409 & new_G2436 & new_G2420 & new_G2472;
  assign new_G2522 = new_G2420 & new_G2454 & new_G2436 & G4526 & new_G2472;
  assign new_G2526 = new_G2454 & new_G2436 & G4526 & new_G2472;
  assign new_G2529 = new_G2454 & G4526 & new_G2472;
  assign new_G2531 = G4526 & new_G2472;
  assign new_G5944 = ~new_G5940;
  assign new_G5952 = ~new_G5948;
  assign new_G5960 = ~new_G5956;
  assign new_G5968 = ~new_G5964;
  assign new_G2555 = ~new_G5972 | ~new_G5975;
  assign new_G5976 = ~new_G5972;
  assign new_G2559 = ~new_G5980 | ~new_G5983;
  assign new_G5984 = ~new_G5980;
  assign new_G2753 = ~new_G2749;
  assign new_G2771 = new_G2643 & new_G2655 & new_G2676 & new_G2742 & new_G2701;
  assign new_G2791 = new_G2701 & new_G2655 & new_G2742 & new_G2676;
  assign new_G2797 = new_G2701 & new_G2742 & new_G2676;
  assign new_G2807 = new_G2742 & new_G2701;
  assign new_G6114 = ~new_G6110;
  assign new_G6172 = ~new_G6168;
  assign new_G6250 = ~new_G6246;
  assign new_G6260 = ~new_G6256;
  assign new_G6346 = ~new_G6342;
  assign new_G6356 = ~new_G6352;
  assign new_G3127 = ~new_G3123;
  assign new_G3156 = new_G3123 & new_G3136;
  assign new_G3259 = new_G3223 | new_G3258;
  assign new_G3466 = new_G3431 & new_G3446;
  assign new_G6646 = ~new_G6642;
  assign new_G6654 = ~new_G6650;
  assign new_G6662 = ~new_G6658;
  assign new_G6670 = ~new_G6666;
  assign new_G3483 = ~new_G6674 | ~new_G6677;
  assign new_G6678 = ~new_G6674;
  assign new_G3487 = ~new_G6682 | ~new_G6685;
  assign new_G6686 = ~new_G6682;
  assign new_G3582 = ~new_G3579;
  assign new_G3586 = ~new_G3583;
  assign new_G3590 = ~new_G3587;
  assign new_G3594 = ~new_G3591;
  assign new_G3597 = ~new_G3595 & ~new_G3596;
  assign new_G3600 = ~new_G3598 & ~new_G3599;
  assign new_G3602 = new_G3579 & new_G3536 & new_G3527;
  assign new_G3605 = new_G3583 & new_G3540 & new_G3531;
  assign new_G3608 = new_G3587 & new_G3559 & new_G3550;
  assign new_G3611 = new_G3591 & new_G3563 & new_G3554;
  assign new_G4023 = ~new_G4020;
  assign new_G6982 = ~new_G6978;
  assign new_G7040 = ~new_G7036;
  assign new_G7118 = ~new_G7114;
  assign new_G7128 = ~new_G7124;
  assign new_G4089 = new_G4004 & new_G4020;
  assign new_G4250 = ~new_G4247;
  assign new_G4254 = ~new_G4251;
  assign new_G4258 = ~new_G4255;
  assign new_G4262 = ~new_G4259;
  assign new_G4272 = new_G4247 & new_G4189 & new_G4180;
  assign new_G4275 = new_G4251 & new_G4193 & new_G4184;
  assign new_G4278 = new_G4255 & new_G4212 & new_G4203;
  assign new_G4281 = new_G4259 & new_G4216 & new_G4207;
  assign new_G4285 = ~new_G4283 & ~new_G4284;
  assign new_G4288 = ~new_G4286 & ~new_G4287;
  assign new_G4360 = ~new_G4356;
  assign new_G4380 = ~new_G4369 | ~G89;
  assign new_G4386 = new_G4356 & new_G4369;
  assign new_G7442 = ~new_G7438;
  assign new_G4609 = ~new_G4606;
  assign new_G4613 = ~new_G4610;
  assign new_G4617 = ~new_G4614;
  assign new_G4621 = ~new_G4618;
  assign new_G4624 = ~new_G4622 & ~new_G4623;
  assign new_G4627 = ~new_G4625 & ~new_G4626;
  assign new_G4629 = new_G4606 & new_G4563 & new_G4554;
  assign new_G4632 = new_G4610 & new_G4567 & new_G4558;
  assign new_G4635 = new_G4614 & new_G4586 & new_G4577;
  assign new_G4638 = new_G4618 & new_G4590 & new_G4581;
  assign new_G4836 = new_G2472;
  assign new_G4949 = ~new_G4947 | ~new_G4948;
  assign new_G4990 = ~new_G4988 | ~new_G4989;
  assign new_G5020 = ~new_G5011 | ~new_G5018;
  assign new_G5108 = ~new_G5099 | ~new_G5106;
  assign new_G5590 = ~new_G5581 | ~new_G5588;
  assign new_G5678 = ~new_G5669 | ~new_G5676;
  assign new_G6084 = ~new_G6080;
  assign new_G6094 = ~new_G6090;
  assign new_G6104 = ~new_G6100;
  assign new_G6142 = ~new_G6138;
  assign new_G6152 = ~new_G6148;
  assign new_G6162 = ~new_G6158;
  assign new_G6206 = new_G2742;
  assign new_G6220 = ~new_G6216;
  assign new_G6230 = ~new_G6226;
  assign new_G6240 = ~new_G6236;
  assign new_G6328 = ~new_G6324;
  assign new_G6294 = new_G2742;
  assign new_G6308 = ~new_G6304;
  assign new_G6318 = ~new_G6314;
  assign new_G6362 = ~new_G6360 | ~new_G6361;
  assign new_G6840 = ~new_G6817 | ~new_G6818;
  assign new_G6848 = ~new_G6827 | ~new_G6828;
  assign new_G6952 = ~new_G6948;
  assign new_G6962 = ~new_G6958;
  assign new_G6972 = ~new_G6968;
  assign new_G7010 = ~new_G7006;
  assign new_G7020 = ~new_G7016;
  assign new_G7030 = ~new_G7026;
  assign new_G7078 = ~new_G7074;
  assign new_G7088 = ~new_G7084;
  assign new_G7098 = ~new_G7094;
  assign new_G7108 = ~new_G7104;
  assign new_G7196 = ~new_G7192;
  assign new_G7166 = ~new_G7162;
  assign new_G7176 = ~new_G7172;
  assign new_G7186 = ~new_G7182;
  assign new_G7448 = ~new_G7446 | ~new_G7447;
  assign new_G7458 = ~new_G7456 | ~new_G7457;
  assign new_G254 = new_G3046 & new_G3249;
  assign new_G260 = new_G3046 & new_G3249;
  assign new_G1987 = ~new_G1985 | ~new_G1986;
  assign new_G1994 = ~new_G1992 | ~new_G1993;
  assign new_G2002 = ~new_G2001;
  assign new_G962 = new_G933 & new_G924;
  assign new_G1751 = new_G1730 & new_G1721;
  assign new_G1990 = ~new_G1988 | ~new_G1989;
  assign new_G1997 = ~new_G1995 | ~new_G1996;
  assign new_G2499 = ~new_G2495;
  assign new_G2536 = new_G2515 & new_G2487;
  assign new_G5943 = ~new_G5937;
  assign new_G2542 = ~new_G5937 | ~new_G5944;
  assign new_G5951 = ~new_G5945;
  assign new_G2545 = ~new_G5945 | ~new_G5952;
  assign new_G5959 = ~new_G5953;
  assign new_G2549 = ~new_G5953 | ~new_G5960;
  assign new_G5967 = ~new_G5961;
  assign new_G2552 = ~new_G5961 | ~new_G5968;
  assign new_G2556 = ~new_G5969 | ~new_G5976;
  assign new_G2560 = ~new_G5977 | ~new_G5984;
  assign new_G2761 = ~new_G2757;
  assign new_G2784 = ~new_G2780;
  assign new_G2853 = new_G2749 & new_G2780;
  assign new_G3135 = ~new_G3131;
  assign new_G3146 = ~new_G3143;
  assign new_G3163 = new_G3123 & new_G3143;
  assign new_G3467 = new_G3453 & new_G3431;
  assign new_G6645 = ~new_G6639;
  assign new_G3470 = ~new_G6639 | ~new_G6646;
  assign new_G6653 = ~new_G6647;
  assign new_G3473 = ~new_G6647 | ~new_G6654;
  assign new_G6661 = ~new_G6655;
  assign new_G3477 = ~new_G6655 | ~new_G6662;
  assign new_G6669 = ~new_G6663;
  assign new_G3480 = ~new_G6663 | ~new_G6670;
  assign new_G3484 = ~new_G6671 | ~new_G6678;
  assign new_G3488 = ~new_G6679 | ~new_G6686;
  assign new_G3601 = new_G3582 & new_G3531 & new_G3536;
  assign new_G3604 = new_G3586 & new_G3527 & new_G3540;
  assign new_G3607 = new_G3590 & new_G3554 & new_G3559;
  assign new_G3610 = new_G3594 & new_G3550 & new_G3563;
  assign new_G4032 = ~new_G4028;
  assign new_G4090 = new_G4004 & new_G4028;
  assign new_G4271 = new_G4250 & new_G4184 & new_G4189;
  assign new_G4274 = new_G4254 & new_G4180 & new_G4193;
  assign new_G4277 = new_G4258 & new_G4207 & new_G4212;
  assign new_G4280 = new_G4262 & new_G4203 & new_G4216;
  assign new_G4368 = ~new_G4364;
  assign new_G4379 = ~new_G4376;
  assign new_G4387 = new_G4356 & new_G4376;
  assign new_G4628 = new_G4609 & new_G4558 & new_G4563;
  assign new_G4631 = new_G4613 & new_G4554 & new_G4567;
  assign new_G4634 = new_G4617 & new_G4581 & new_G4586;
  assign new_G4637 = new_G4621 & new_G4577 & new_G4590;
  assign new_G4841 = new_G2522 | new_G2520 | new_G2519 | new_G2431 | new_G2518;
  assign new_G4849 = new_G2526 | new_G2524 | new_G2448 | new_G2523;
  assign new_G4857 = new_G2529 | new_G2465 | new_G2527;
  assign new_G4865 = new_G2481 | new_G2531;
  assign new_G5021 = ~new_G5019 | ~new_G5020;
  assign new_G5028 = ~new_G5024;
  assign new_G5109 = ~new_G5107 | ~new_G5108;
  assign new_G5116 = ~new_G5112;
  assign new_G5369 = ~new_G1313 | ~new_G1310;
  assign new_G5377 = ~new_G1319 | ~new_G1316;
  assign new_G5385 = ~new_G1325 | ~new_G1322;
  assign new_G5472 = ~new_G5468;
  assign new_G5473 = ~new_G5468 | ~new_G5471;
  assign new_G5530 = ~new_G5526;
  assign new_G5531 = ~new_G5526 | ~new_G5529;
  assign new_G5591 = ~new_G5589 | ~new_G5590;
  assign new_G5598 = ~new_G5594;
  assign new_G5679 = ~new_G5677 | ~new_G5678;
  assign new_G5686 = ~new_G5682;
  assign new_G6060 = new_G2768 | new_G2804;
  assign new_G6074 = ~new_G6070;
  assign new_G6118 = ~new_G2768;
  assign new_G6132 = ~new_G6128;
  assign new_G6176 = new_G2797 | new_G2796 | new_G2693 | new_G2795;
  assign new_G6186 = new_G2801 | new_G2807;
  assign new_G6196 = new_G2791 | new_G2790 | new_G2789 | new_G2670 | new_G2788;
  assign new_G6268 = ~new_G6264;
  assign new_G6269 = ~new_G6264 | ~new_G6267;
  assign new_G6274 = ~new_G2801;
  assign new_G6288 = ~new_G6284;
  assign new_G6337 = ~new_G4288 | ~new_G4285;
  assign new_G6829 = ~new_G3600 | ~new_G3597;
  assign new_G6928 = new_G4017 | new_G4051;
  assign new_G6942 = ~new_G6938;
  assign new_G6986 = ~new_G4017;
  assign new_G7000 = ~new_G6996;
  assign new_G7048 = ~new_G7044;
  assign new_G7049 = ~new_G7044 | ~new_G7047;
  assign new_G7054 = new_G4048 | new_G4052;
  assign new_G7068 = ~new_G7064;
  assign new_G7136 = ~new_G7132;
  assign new_G7137 = ~new_G7132 | ~new_G7135;
  assign new_G7142 = ~new_G4048;
  assign new_G7156 = ~new_G7152;
  assign new_G7433 = ~new_G4627 | ~new_G4624;
  assign new_G242 = new_G1982 & new_G1146;
  assign new_G3151 = ~new_G3135 | ~new_G3127;
  assign new_G257 = new_G3249 & new_G3035 & new_G3156 & G89 & new_G4386;
  assign new_G263 = new_G3249 & new_G3035 & new_G3156 & G89 & new_G4386;
  assign new_G266 = new_G1790 & new_G997;
  assign new_G1991 = ~new_G1990;
  assign new_G1998 = ~new_G1997;
  assign new_G3489 = ~new_G3487 | ~new_G3488;
  assign new_G371 = ~new_G4836 | ~new_G4839;
  assign new_G4840 = ~new_G4836;
  assign new_G2561 = ~new_G2559 | ~new_G2560;
  assign new_G2532 = new_G2487 & new_G2508;
  assign new_G2537 = new_G2495 | new_G2536;
  assign new_G2541 = ~new_G5940 | ~new_G5943;
  assign new_G2544 = ~new_G5948 | ~new_G5951;
  assign new_G2548 = ~new_G5956 | ~new_G5959;
  assign new_G2551 = ~new_G5964 | ~new_G5967;
  assign new_G2557 = ~new_G2555 | ~new_G2556;
  assign new_G2563 = new_G2508 & G4526;
  assign new_G2577 = ~new_G2499 | ~new_G2491;
  assign new_G2775 = ~new_G2771;
  assign new_G2806 = ~new_G2771 | ~G4526;
  assign new_G2808 = ~new_G2761 | ~new_G2753;
  assign new_G2852 = new_G2749 & new_G2771;
  assign new_G2854 = new_G2757 | new_G2853;
  assign new_G6366 = ~new_G6362;
  assign new_G4381 = ~new_G4368 | ~new_G4360;
  assign new_G3164 = new_G3131 | new_G3163;
  assign new_G3241 = new_G3035 & new_G3156 & G89 & new_G4386;
  assign new_G3468 = new_G3437 | new_G3467;
  assign new_G3469 = ~new_G6642 | ~new_G6645;
  assign new_G3472 = ~new_G6650 | ~new_G6653;
  assign new_G3476 = ~new_G6658 | ~new_G6661;
  assign new_G3479 = ~new_G6666 | ~new_G6669;
  assign new_G3485 = ~new_G3483 | ~new_G3484;
  assign new_G3603 = ~new_G3601 & ~new_G3602;
  assign new_G3606 = ~new_G3604 & ~new_G3605;
  assign new_G3609 = ~new_G3607 & ~new_G3608;
  assign new_G3612 = ~new_G3610 & ~new_G3611;
  assign new_G6844 = ~new_G6840;
  assign new_G6852 = ~new_G6848;
  assign new_G4091 = new_G4010 | new_G4090;
  assign new_G4273 = ~new_G4271 & ~new_G4272;
  assign new_G4276 = ~new_G4274 & ~new_G4275;
  assign new_G4279 = ~new_G4277 & ~new_G4278;
  assign new_G4282 = ~new_G4280 & ~new_G4281;
  assign new_G4382 = new_G4379 & new_G4380;
  assign new_G4388 = new_G4364 | new_G4387;
  assign new_G7452 = ~new_G7448;
  assign new_G7462 = ~new_G7458;
  assign new_G4630 = ~new_G4628 & ~new_G4629;
  assign new_G4633 = ~new_G4631 & ~new_G4632;
  assign new_G4636 = ~new_G4634 & ~new_G4635;
  assign new_G4639 = ~new_G4637 & ~new_G4638;
  assign new_G4955 = ~new_G4949;
  assign new_G4958 = ~new_G4949 | ~new_G4956;
  assign new_G4996 = ~new_G4990;
  assign new_G4999 = ~new_G4990 | ~new_G4997;
  assign new_G5474 = ~new_G5465 | ~new_G5472;
  assign new_G5532 = ~new_G5523 | ~new_G5530;
  assign new_G6210 = ~new_G6206;
  assign new_G6270 = ~new_G6261 | ~new_G6268;
  assign new_G6298 = ~new_G6294;
  assign new_G7050 = ~new_G7041 | ~new_G7048;
  assign new_G7138 = ~new_G7129 | ~new_G7136;
  assign new_G3471 = ~new_G3469 | ~new_G3470;
  assign new_G3478 = ~new_G3476 | ~new_G3477;
  assign new_G3486 = ~new_G3485;
  assign new_G372 = ~new_G4833 | ~new_G4840;
  assign new_G2543 = ~new_G2541 | ~new_G2542;
  assign new_G2550 = ~new_G2548 | ~new_G2549;
  assign new_G2558 = ~new_G2557;
  assign new_G4847 = ~new_G4841;
  assign new_G387 = ~new_G4841 | ~new_G4848;
  assign new_G4855 = ~new_G4849;
  assign new_G390 = ~new_G4849 | ~new_G4856;
  assign new_G4863 = ~new_G4857;
  assign new_G393 = ~new_G4857 | ~new_G4864;
  assign new_G4871 = ~new_G4865;
  assign new_G396 = ~new_G4865 | ~new_G4872;
  assign new_G965 = ~new_G962;
  assign new_G5375 = ~new_G5369;
  assign new_G1327 = ~new_G5369 | ~new_G5376;
  assign new_G5383 = ~new_G5377;
  assign new_G1330 = ~new_G5377 | ~new_G5384;
  assign new_G5391 = ~new_G5385;
  assign new_G1333 = ~new_G5385 | ~new_G5392;
  assign new_G1754 = ~new_G1751;
  assign new_G2546 = ~new_G2544 | ~new_G2545;
  assign new_G2553 = ~new_G2551 | ~new_G2552;
  assign new_G2564 = new_G2515 | new_G2563;
  assign new_G2809 = new_G2784 & new_G2806;
  assign new_G2813 = new_G2784 & new_G2775;
  assign new_G6345 = ~new_G6337;
  assign new_G2860 = ~new_G6337 | ~new_G6346;
  assign new_G3474 = ~new_G3472 | ~new_G3473;
  assign new_G3481 = ~new_G3479 | ~new_G3480;
  assign new_G6835 = ~new_G6829;
  assign new_G3614 = ~new_G6829 | ~new_G6836;
  assign new_G4053 = new_G4032 & new_G4023;
  assign new_G7441 = ~new_G7433;
  assign new_G4516 = ~new_G7433 | ~new_G7442;
  assign new_G4957 = ~new_G4952 | ~new_G4955;
  assign new_G4998 = ~new_G4993 | ~new_G4996;
  assign new_G5027 = ~new_G5021;
  assign new_G5030 = ~new_G5021 | ~new_G5028;
  assign new_G5115 = ~new_G5109;
  assign new_G5118 = ~new_G5109 | ~new_G5116;
  assign new_G5475 = ~new_G5473 | ~new_G5474;
  assign new_G5533 = ~new_G5531 | ~new_G5532;
  assign new_G5597 = ~new_G5591;
  assign new_G5600 = ~new_G5591 | ~new_G5598;
  assign new_G5685 = ~new_G5679;
  assign new_G5688 = ~new_G5679 | ~new_G5686;
  assign new_G6064 = ~new_G6060;
  assign new_G6065 = ~new_G6060 | ~new_G6063;
  assign new_G6122 = ~new_G6118;
  assign new_G6123 = ~new_G6118 | ~new_G6121;
  assign new_G6180 = ~new_G6176;
  assign new_G6181 = ~new_G6176 | ~new_G6179;
  assign new_G6190 = ~new_G6186;
  assign new_G6200 = ~new_G6196;
  assign new_G6271 = ~new_G6269 | ~new_G6270;
  assign new_G6278 = ~new_G6274;
  assign new_G6347 = ~new_G4276 | ~new_G4273;
  assign new_G6357 = ~new_G4282 | ~new_G4279;
  assign new_G6837 = ~new_G3606 | ~new_G3603;
  assign new_G6845 = ~new_G3612 | ~new_G3609;
  assign new_G6932 = ~new_G6928;
  assign new_G6933 = ~new_G6928 | ~new_G6931;
  assign new_G6990 = ~new_G6986;
  assign new_G6991 = ~new_G6986 | ~new_G6989;
  assign new_G7051 = ~new_G7049 | ~new_G7050;
  assign new_G7058 = ~new_G7054;
  assign new_G7139 = ~new_G7137 | ~new_G7138;
  assign new_G7146 = ~new_G7142;
  assign new_G7443 = ~new_G4639 | ~new_G4636;
  assign new_G7453 = ~new_G4633 | ~new_G4630;
  assign new_G243 = new_G1146 & new_G3468 & new_G1974;
  assign new_G244 = new_G1146 & new_G1974 & new_G2537 & new_G3466;
  assign new_G245 = new_G1146 & new_G1974 & new_G3466 & G4526 & new_G2532;
  assign new_G255 = new_G3249 & new_G3164 & new_G3035;
  assign new_G256 = new_G3249 & new_G3035 & new_G4388 & new_G3156;
  assign new_G261 = new_G3249 & new_G3164 & new_G3035;
  assign new_G262 = new_G3249 & new_G3035 & new_G4388 & new_G3156;
  assign new_G267 = new_G997 & new_G4091 & new_G1788;
  assign new_G268 = new_G997 & new_G1788 & new_G2854 & new_G4089;
  assign new_G269 = new_G997 & new_G1788 & new_G4089 & G4526 & new_G2852;
  assign new_G3475 = ~new_G3474;
  assign new_G3482 = ~new_G3481;
  assign G373 = ~new_G371 | ~new_G372;
  assign new_G2547 = ~new_G2546;
  assign new_G2554 = ~new_G2553;
  assign new_G386 = ~new_G4844 | ~new_G4847;
  assign new_G389 = ~new_G4852 | ~new_G4855;
  assign new_G392 = ~new_G4860 | ~new_G4863;
  assign new_G395 = ~new_G4868 | ~new_G4871;
  assign new_G1326 = ~new_G5372 | ~new_G5375;
  assign new_G1329 = ~new_G5380 | ~new_G5383;
  assign new_G1332 = ~new_G5388 | ~new_G5391;
  assign new_G1436 = new_G4091 & new_G1788;
  assign new_G1440 = new_G1788 & new_G2854 & new_G4089;
  assign new_G1445 = new_G1788 & new_G4089 & G4526 & new_G2852;
  assign new_G1450 = new_G2854 & new_G4089;
  assign new_G1454 = new_G4089 & G4526 & new_G2852;
  assign new_G2859 = ~new_G6342 | ~new_G6345;
  assign new_G4385 = ~new_G4382;
  assign new_G3148 = new_G4382 & new_G4364;
  assign new_G3239 = new_G3164 & new_G3035;
  assign new_G3240 = new_G3035 & new_G4388 & new_G3156;
  assign new_G3265 = new_G3468 & new_G1974;
  assign new_G3267 = new_G1974 & new_G2537 & new_G3466;
  assign new_G3270 = new_G1974 & new_G3466 & G4526 & new_G2532;
  assign new_G3274 = new_G2537 & new_G3466;
  assign new_G3277 = new_G3466 & G4526 & new_G2532;
  assign new_G3613 = ~new_G6832 | ~new_G6835;
  assign new_G4515 = ~new_G7438 | ~new_G7441;
  assign new_G4959 = ~new_G4957 | ~new_G4958;
  assign new_G5000 = ~new_G4998 | ~new_G4999;
  assign new_G5029 = ~new_G5024 | ~new_G5027;
  assign new_G5117 = ~new_G5112 | ~new_G5115;
  assign new_G5599 = ~new_G5594 | ~new_G5597;
  assign new_G5687 = ~new_G5682 | ~new_G5685;
  assign new_G6066 = ~new_G6057 | ~new_G6064;
  assign new_G6124 = ~new_G6115 | ~new_G6122;
  assign new_G6182 = ~new_G6173 | ~new_G6180;
  assign new_G6934 = ~new_G6925 | ~new_G6932;
  assign new_G6992 = ~new_G6983 | ~new_G6990;
  assign G246 = new_G245 | new_G244 | new_G243 | new_G241 | new_G242;
  assign G258 = new_G257 | new_G256 | new_G255 | new_G3259 | new_G254;
  assign G264 = new_G263 | new_G262 | new_G261 | new_G3259 | new_G260;
  assign G270 = new_G269 | new_G268 | new_G267 | new_G265 | new_G266;
  assign new_G375 = new_G2564 & new_G2543;
  assign new_G378 = new_G2564 & new_G2550;
  assign new_G381 = new_G2564 & new_G2558;
  assign new_G384 = new_G2564 & new_G2406;
  assign G388 = ~new_G386 | ~new_G387;
  assign G391 = ~new_G389 | ~new_G390;
  assign G394 = ~new_G392 | ~new_G393;
  assign G397 = ~new_G395 | ~new_G396;
  assign new_G1328 = ~new_G1326 | ~new_G1327;
  assign new_G1331 = ~new_G1329 | ~new_G1330;
  assign new_G1334 = ~new_G1332 | ~new_G1333;
  assign new_G1447 = new_G1445 | new_G1440 | new_G1790 | new_G1436;
  assign new_G1766 = new_G1454 | new_G4091 | new_G1450;
  assign new_G2571 = ~new_G2564;
  assign new_G2579 = new_G2577 & new_G2564;
  assign new_G2812 = ~new_G2809;
  assign new_G2816 = ~new_G2813;
  assign new_G2851 = new_G2809 & new_G2757;
  assign new_G2861 = ~new_G2859 | ~new_G2860;
  assign new_G6355 = ~new_G6347;
  assign new_G2863 = ~new_G6347 | ~new_G6356;
  assign new_G6365 = ~new_G6357;
  assign new_G2866 = ~new_G6357 | ~new_G6366;
  assign new_G3147 = new_G4381 & new_G4385;
  assign new_G3242 = new_G3241 | new_G3240 | new_G3046 | new_G3239;
  assign new_G3271 = new_G3270 | new_G3267 | new_G1982 | new_G3265;
  assign new_G3279 = new_G3277 | new_G3468 | new_G3274;
  assign new_G3615 = ~new_G3613 | ~new_G3614;
  assign new_G6843 = ~new_G6837;
  assign new_G3617 = ~new_G6837 | ~new_G6844;
  assign new_G6851 = ~new_G6845;
  assign new_G3620 = ~new_G6845 | ~new_G6852;
  assign new_G4056 = ~new_G4053;
  assign new_G4517 = ~new_G4515 | ~new_G4516;
  assign new_G7451 = ~new_G7443;
  assign new_G4519 = ~new_G7443 | ~new_G7452;
  assign new_G7461 = ~new_G7453;
  assign new_G4522 = ~new_G7453 | ~new_G7462;
  assign new_G5031 = ~new_G5029 | ~new_G5030;
  assign new_G5119 = ~new_G5117 | ~new_G5118;
  assign new_G5481 = ~new_G5475;
  assign new_G5484 = ~new_G5475 | ~new_G5482;
  assign new_G5539 = ~new_G5533;
  assign new_G5542 = ~new_G5533 | ~new_G5540;
  assign new_G5601 = ~new_G5599 | ~new_G5600;
  assign new_G5689 = ~new_G5687 | ~new_G5688;
  assign new_G6067 = ~new_G6065 | ~new_G6066;
  assign new_G6125 = ~new_G6123 | ~new_G6124;
  assign new_G6183 = ~new_G6181 | ~new_G6182;
  assign new_G6277 = ~new_G6271;
  assign new_G6280 = ~new_G6271 | ~new_G6278;
  assign new_G6935 = ~new_G6933 | ~new_G6934;
  assign new_G6993 = ~new_G6991 | ~new_G6992;
  assign new_G7057 = ~new_G7051;
  assign new_G7060 = ~new_G7051 | ~new_G7058;
  assign new_G7145 = ~new_G7139;
  assign new_G7148 = ~new_G7139 | ~new_G7146;
  assign new_G4968 = ~new_G4959 | ~new_G4966;
  assign new_G5009 = ~new_G5000 | ~new_G5007;
  assign new_G2850 = new_G2808 & new_G2812;
  assign new_G2862 = ~new_G6352 | ~new_G6355;
  assign new_G2865 = ~new_G6362 | ~new_G6365;
  assign new_G3149 = new_G3147 | new_G3148;
  assign new_G3243 = ~new_G3228 | ~new_G3242;
  assign new_G3616 = ~new_G6840 | ~new_G6843;
  assign new_G3619 = ~new_G6848 | ~new_G6851;
  assign new_G4518 = ~new_G7448 | ~new_G7451;
  assign new_G4521 = ~new_G7458 | ~new_G7461;
  assign new_G4965 = ~new_G4959;
  assign new_G5006 = ~new_G5000;
  assign new_G5483 = ~new_G5478 | ~new_G5481;
  assign new_G5541 = ~new_G5536 | ~new_G5539;
  assign new_G6279 = ~new_G6274 | ~new_G6277;
  assign new_G7059 = ~new_G7054 | ~new_G7057;
  assign new_G7147 = ~new_G7142 | ~new_G7145;
  assign new_G374 = new_G2547 & new_G2571;
  assign new_G377 = new_G2554 & new_G2571;
  assign new_G380 = new_G2561 & new_G2571;
  assign new_G383 = new_G2400 & new_G2571;
  assign new_G955 = ~new_G920 | ~new_G1447;
  assign new_G4967 = ~new_G4962 | ~new_G4965;
  assign new_G5008 = ~new_G5003 | ~new_G5006;
  assign new_G975 = new_G1447;
  assign new_G1136 = new_G1038 & new_G1074 & new_G1055 & new_G3271 & new_G1093;
  assign new_G1140 = new_G1074 & new_G1055 & new_G3271 & new_G1093;
  assign new_G1143 = new_G1074 & new_G3271 & new_G1093;
  assign new_G1145 = new_G3271 & new_G1093;
  assign new_G1160 = new_G1122 & new_G3271;
  assign new_G1771 = ~new_G1766;
  assign new_G1964 = new_G1869 & new_G1903 & new_G1885 & new_G3279 & new_G1921;
  assign new_G1968 = new_G1903 & new_G1885 & new_G3279 & new_G1921;
  assign new_G1971 = new_G1903 & new_G3279 & new_G1921;
  assign new_G1973 = new_G3279 & new_G1921;
  assign new_G2007 = new_G1950 & new_G3279;
  assign new_G2578 = new_G2495 & new_G2571;
  assign new_G2864 = ~new_G2862 | ~new_G2863;
  assign new_G2867 = ~new_G2865 | ~new_G2866;
  assign new_G3150 = ~new_G3136 | ~new_G3149;
  assign new_G3245 = new_G3238 & new_G3243;
  assign new_G3618 = ~new_G3616 | ~new_G3617;
  assign new_G3621 = ~new_G3619 | ~new_G3620;
  assign new_G4067 = new_G2850 | new_G2851;
  assign new_G4520 = ~new_G4518 | ~new_G4519;
  assign new_G4523 = ~new_G4521 | ~new_G4522;
  assign new_G4713 = new_G3279;
  assign new_G4753 = new_G3271;
  assign new_G5037 = ~new_G5031;
  assign new_G5040 = ~new_G5031 | ~new_G5038;
  assign new_G5125 = ~new_G5119;
  assign new_G5128 = ~new_G5119 | ~new_G5126;
  assign new_G5485 = ~new_G5483 | ~new_G5484;
  assign new_G5543 = ~new_G5541 | ~new_G5542;
  assign new_G5607 = ~new_G5601;
  assign new_G5610 = ~new_G5601 | ~new_G5608;
  assign new_G5695 = ~new_G5689;
  assign new_G5698 = ~new_G5689 | ~new_G5696;
  assign new_G6073 = ~new_G6067;
  assign new_G6076 = ~new_G6067 | ~new_G6074;
  assign new_G6131 = ~new_G6125;
  assign new_G6134 = ~new_G6125 | ~new_G6132;
  assign new_G6189 = ~new_G6183;
  assign new_G6192 = ~new_G6183 | ~new_G6190;
  assign new_G6281 = ~new_G6279 | ~new_G6280;
  assign new_G6941 = ~new_G6935;
  assign new_G6944 = ~new_G6935 | ~new_G6942;
  assign new_G6999 = ~new_G6993;
  assign new_G7002 = ~new_G6993 | ~new_G7000;
  assign new_G7061 = ~new_G7059 | ~new_G7060;
  assign new_G7149 = ~new_G7147 | ~new_G7148;
  assign G376 = new_G374 | new_G375;
  assign G379 = new_G377 | new_G378;
  assign G382 = new_G380 | new_G381;
  assign G385 = new_G383 | new_G384;
  assign new_G958 = new_G933 & new_G955;
  assign new_G967 = ~new_G4967 | ~new_G4968;
  assign new_G971 = ~new_G5008 | ~new_G5009;
  assign new_G1161 = new_G1129 | new_G1160;
  assign new_G2008 = new_G1957 | new_G2007;
  assign new_G2580 = new_G2578 | new_G2579;
  assign new_G2868 = new_G2867 & new_G2864 & new_G1331 & new_G2861;
  assign new_G3152 = new_G3146 & new_G3150;
  assign new_G4443 = new_G3621 & new_G3618 & new_G1328 & new_G1334;
  assign new_G4524 = new_G4523 & new_G4520 & new_G3615 & new_G4517;
  assign new_G4721 = new_G1964 | new_G1962 | new_G1961 | new_G1880 | new_G1960;
  assign new_G4729 = new_G1968 | new_G1966 | new_G1897 | new_G1965;
  assign new_G4737 = new_G1971 | new_G1914 | new_G1969;
  assign new_G4745 = new_G1929 | new_G1973;
  assign new_G4761 = new_G1136 | new_G1134 | new_G1133 | new_G1050 | new_G1132;
  assign new_G4769 = new_G1140 | new_G1138 | new_G1068 | new_G1137;
  assign new_G4777 = new_G1143 | new_G1086 | new_G1141;
  assign new_G4785 = new_G1102 | new_G1145;
  assign new_G5039 = ~new_G5034 | ~new_G5037;
  assign new_G5127 = ~new_G5122 | ~new_G5125;
  assign new_G5609 = ~new_G5604 | ~new_G5607;
  assign new_G5697 = ~new_G5692 | ~new_G5695;
  assign new_G6075 = ~new_G6070 | ~new_G6073;
  assign new_G6133 = ~new_G6128 | ~new_G6131;
  assign new_G6191 = ~new_G6186 | ~new_G6189;
  assign new_G6943 = ~new_G6938 | ~new_G6941;
  assign new_G7001 = ~new_G6996 | ~new_G6999;
  assign new_G3248 = ~new_G3245;
  assign new_G248 = new_G3245 & new_G3223;
  assign new_G4719 = ~new_G4713;
  assign new_G294 = ~new_G4713 | ~new_G4720;
  assign new_G4759 = ~new_G4753;
  assign new_G323 = ~new_G4753 | ~new_G4760;
  assign new_G980 = ~new_G975;
  assign new_G4072 = ~new_G4067;
  assign new_G5041 = ~new_G5039 | ~new_G5040;
  assign new_G5129 = ~new_G5127 | ~new_G5128;
  assign new_G5491 = ~new_G5485;
  assign new_G5494 = ~new_G5485 | ~new_G5492;
  assign new_G5549 = ~new_G5543;
  assign new_G5552 = ~new_G5543 | ~new_G5550;
  assign new_G5611 = ~new_G5609 | ~new_G5610;
  assign new_G5699 = ~new_G5697 | ~new_G5698;
  assign new_G6077 = ~new_G6075 | ~new_G6076;
  assign new_G6135 = ~new_G6133 | ~new_G6134;
  assign new_G6193 = ~new_G6191 | ~new_G6192;
  assign new_G6287 = ~new_G6281;
  assign new_G6290 = ~new_G6281 | ~new_G6288;
  assign new_G6945 = ~new_G6943 | ~new_G6944;
  assign new_G7003 = ~new_G7001 | ~new_G7002;
  assign new_G7067 = ~new_G7061;
  assign new_G7070 = ~new_G7061 | ~new_G7068;
  assign new_G7155 = ~new_G7149;
  assign new_G7158 = ~new_G7149 | ~new_G7156;
  assign new_G247 = new_G3244 & new_G3248;
  assign new_G3155 = ~new_G3152;
  assign new_G251 = new_G3152 & new_G3131;
  assign new_G272 = new_G1176 & new_G1161;
  assign new_G961 = ~new_G958;
  assign new_G275 = new_G958 & new_G908;
  assign new_G293 = ~new_G4716 | ~new_G4719;
  assign new_G297 = new_G2008 & new_G1987;
  assign new_G300 = new_G2008 & new_G1994;
  assign new_G303 = new_G2008 & new_G2002;
  assign new_G306 = new_G2008 & new_G1856;
  assign new_G4727 = ~new_G4721;
  assign new_G309 = ~new_G4721 | ~new_G4728;
  assign new_G4735 = ~new_G4729;
  assign new_G312 = ~new_G4729 | ~new_G4736;
  assign new_G4743 = ~new_G4737;
  assign new_G315 = ~new_G4737 | ~new_G4744;
  assign new_G4751 = ~new_G4745;
  assign new_G318 = ~new_G4745 | ~new_G4752;
  assign new_G322 = ~new_G4756 | ~new_G4759;
  assign new_G4767 = ~new_G4761;
  assign new_G326 = ~new_G4761 | ~new_G4768;
  assign new_G4775 = ~new_G4769;
  assign new_G329 = ~new_G4769 | ~new_G4776;
  assign new_G4783 = ~new_G4777;
  assign new_G332 = ~new_G4777 | ~new_G4784;
  assign new_G4791 = ~new_G4785;
  assign new_G335 = ~new_G4785 | ~new_G4792;
  assign G412 = ~new_G4443;
  assign G414 = ~new_G4524;
  assign G416 = ~new_G2868;
  assign new_G2881 = new_G2868 & new_G4443 & new_G4524;
  assign new_G993 = new_G975 & new_G971 & new_G962;
  assign new_G994 = new_G975 & new_G967 & new_G965;
  assign new_G1166 = ~new_G1161;
  assign new_G1171 = new_G1161 & new_G1155;
  assign new_G1174 = new_G1161 & new_G1023;
  assign new_G2014 = ~new_G2008;
  assign new_G3459 = new_G3365 & new_G3399 & new_G3381 & new_G2580 & new_G3417;
  assign new_G3462 = new_G3399 & new_G3381 & new_G2580 & new_G3417;
  assign new_G3464 = new_G3399 & new_G2580 & new_G3417;
  assign new_G3465 = new_G2580 & new_G3417;
  assign new_G3490 = new_G3446 & new_G2580;
  assign new_G4793 = new_G2580;
  assign new_G5493 = ~new_G5488 | ~new_G5491;
  assign new_G5551 = ~new_G5546 | ~new_G5549;
  assign new_G6289 = ~new_G6284 | ~new_G6287;
  assign new_G7069 = ~new_G7064 | ~new_G7067;
  assign new_G7157 = ~new_G7152 | ~new_G7155;
  assign G249 = new_G247 | new_G248;
  assign new_G250 = new_G3151 & new_G3155;
  assign new_G274 = new_G957 & new_G961;
  assign G295 = ~new_G293 | ~new_G294;
  assign new_G308 = ~new_G4724 | ~new_G4727;
  assign new_G311 = ~new_G4732 | ~new_G4735;
  assign new_G314 = ~new_G4740 | ~new_G4743;
  assign new_G317 = ~new_G4748 | ~new_G4751;
  assign G324 = ~new_G322 | ~new_G323;
  assign new_G325 = ~new_G4764 | ~new_G4767;
  assign new_G328 = ~new_G4772 | ~new_G4775;
  assign new_G331 = ~new_G4780 | ~new_G4783;
  assign new_G334 = ~new_G4788 | ~new_G4791;
  assign new_G417 = new_G2881 & new_G2876 & new_G2878;
  assign new_G991 = new_G980 & new_G971 & new_G933;
  assign new_G992 = new_G980 & new_G967 & new_G929;
  assign new_G3491 = new_G3453 | new_G3490;
  assign new_G4801 = new_G3459 | new_G3458 | new_G3457 | new_G3376 | new_G3456;
  assign new_G4809 = new_G3462 | new_G3461 | new_G3393 | new_G3460;
  assign new_G4817 = new_G3464 | new_G3410 | new_G3463;
  assign new_G4825 = new_G3425 | new_G3465;
  assign new_G5047 = ~new_G5041;
  assign new_G5050 = ~new_G5041 | ~new_G5048;
  assign new_G5135 = ~new_G5129;
  assign new_G5138 = ~new_G5129 | ~new_G5136;
  assign new_G5495 = ~new_G5493 | ~new_G5494;
  assign new_G5553 = ~new_G5551 | ~new_G5552;
  assign new_G5617 = ~new_G5611;
  assign new_G5620 = ~new_G5611 | ~new_G5618;
  assign new_G5705 = ~new_G5699;
  assign new_G5708 = ~new_G5699 | ~new_G5706;
  assign new_G6083 = ~new_G6077;
  assign new_G6086 = ~new_G6077 | ~new_G6084;
  assign new_G6141 = ~new_G6135;
  assign new_G6144 = ~new_G6135 | ~new_G6142;
  assign new_G6199 = ~new_G6193;
  assign new_G6202 = ~new_G6193 | ~new_G6200;
  assign new_G6291 = ~new_G6289 | ~new_G6290;
  assign new_G6951 = ~new_G6945;
  assign new_G6954 = ~new_G6945 | ~new_G6952;
  assign new_G7009 = ~new_G7003;
  assign new_G7012 = ~new_G7003 | ~new_G7010;
  assign new_G7071 = ~new_G7069 | ~new_G7070;
  assign new_G7159 = ~new_G7157 | ~new_G7158;
  assign G252 = new_G250 | new_G251;
  assign new_G271 = new_G1117 & new_G1166;
  assign G276 = new_G274 | new_G275;
  assign new_G296 = new_G1991 & new_G2014;
  assign new_G299 = new_G1998 & new_G2014;
  assign new_G302 = new_G2005 & new_G2014;
  assign new_G305 = new_G1850 & new_G2014;
  assign G310 = ~new_G308 | ~new_G309;
  assign G313 = ~new_G311 | ~new_G312;
  assign G316 = ~new_G314 | ~new_G315;
  assign G319 = ~new_G317 | ~new_G318;
  assign G327 = ~new_G325 | ~new_G326;
  assign G330 = ~new_G328 | ~new_G329;
  assign G333 = ~new_G331 | ~new_G332;
  assign G336 = ~new_G334 | ~new_G335;
  assign new_G4799 = ~new_G4793;
  assign new_G343 = ~new_G4793 | ~new_G4800;
  assign G418 = ~new_G417;
  assign new_G1170 = new_G1158 & new_G1166;
  assign new_G1173 = new_G1019 & new_G1166;
  assign new_G5049 = ~new_G5044 | ~new_G5047;
  assign new_G5137 = ~new_G5132 | ~new_G5135;
  assign new_G5167 = new_G994 | new_G993 | new_G991 | new_G992;
  assign new_G5619 = ~new_G5614 | ~new_G5617;
  assign new_G5707 = ~new_G5702 | ~new_G5705;
  assign new_G6085 = ~new_G6080 | ~new_G6083;
  assign new_G6143 = ~new_G6138 | ~new_G6141;
  assign new_G6201 = ~new_G6196 | ~new_G6199;
  assign new_G6953 = ~new_G6948 | ~new_G6951;
  assign new_G7011 = ~new_G7006 | ~new_G7009;
  assign G273 = new_G271 | new_G272;
  assign G298 = new_G296 | new_G297;
  assign G301 = new_G299 | new_G300;
  assign G304 = new_G302 | new_G303;
  assign G307 = new_G305 | new_G306;
  assign new_G342 = ~new_G4796 | ~new_G4799;
  assign new_G346 = new_G3491 & new_G3471;
  assign new_G349 = new_G3491 & new_G3478;
  assign new_G352 = new_G3491 & new_G3486;
  assign new_G355 = new_G3491 & new_G3350;
  assign new_G4807 = ~new_G4801;
  assign new_G358 = ~new_G4801 | ~new_G4808;
  assign new_G4815 = ~new_G4809;
  assign new_G361 = ~new_G4809 | ~new_G4816;
  assign new_G4823 = ~new_G4817;
  assign new_G364 = ~new_G4817 | ~new_G4824;
  assign new_G4831 = ~new_G4825;
  assign new_G367 = ~new_G4825 | ~new_G4832;
  assign new_G1172 = new_G1170 | new_G1171;
  assign new_G1175 = new_G1173 | new_G1174;
  assign new_G3497 = ~new_G3491;
  assign new_G5051 = ~new_G5049 | ~new_G5050;
  assign new_G5139 = ~new_G5137 | ~new_G5138;
  assign new_G5501 = ~new_G5495;
  assign new_G5504 = ~new_G5495 | ~new_G5502;
  assign new_G5559 = ~new_G5553;
  assign new_G5562 = ~new_G5553 | ~new_G5560;
  assign new_G5621 = ~new_G5619 | ~new_G5620;
  assign new_G5709 = ~new_G5707 | ~new_G5708;
  assign new_G6087 = ~new_G6085 | ~new_G6086;
  assign new_G6145 = ~new_G6143 | ~new_G6144;
  assign new_G6203 = ~new_G6201 | ~new_G6202;
  assign new_G6297 = ~new_G6291;
  assign new_G6300 = ~new_G6291 | ~new_G6298;
  assign new_G6955 = ~new_G6953 | ~new_G6954;
  assign new_G7013 = ~new_G7011 | ~new_G7012;
  assign new_G7077 = ~new_G7071;
  assign new_G7080 = ~new_G7071 | ~new_G7078;
  assign new_G7165 = ~new_G7159;
  assign new_G7168 = ~new_G7159 | ~new_G7166;
  assign G344 = ~new_G342 | ~new_G343;
  assign new_G357 = ~new_G4804 | ~new_G4807;
  assign new_G360 = ~new_G4812 | ~new_G4815;
  assign new_G363 = ~new_G4820 | ~new_G4823;
  assign new_G366 = ~new_G4828 | ~new_G4831;
  assign new_G5173 = ~new_G5167;
  assign G422 = new_G1172;
  assign G469 = new_G1172;
  assign G419 = new_G1175;
  assign G471 = new_G1175;
  assign new_G5503 = ~new_G5498 | ~new_G5501;
  assign new_G5561 = ~new_G5556 | ~new_G5559;
  assign new_G6299 = ~new_G6294 | ~new_G6297;
  assign new_G7079 = ~new_G7074 | ~new_G7077;
  assign new_G7167 = ~new_G7162 | ~new_G7165;
  assign new_G345 = new_G3475 & new_G3497;
  assign new_G348 = new_G3482 & new_G3497;
  assign new_G351 = new_G3489 & new_G3497;
  assign new_G354 = new_G3344 & new_G3497;
  assign G359 = ~new_G357 | ~new_G358;
  assign G362 = ~new_G360 | ~new_G361;
  assign G365 = ~new_G363 | ~new_G364;
  assign G368 = ~new_G366 | ~new_G367;
  assign new_G5057 = ~new_G5051;
  assign new_G5060 = ~new_G5051 | ~new_G5058;
  assign new_G5145 = ~new_G5139;
  assign new_G5148 = ~new_G5139 | ~new_G5146;
  assign new_G5505 = ~new_G5503 | ~new_G5504;
  assign new_G5563 = ~new_G5561 | ~new_G5562;
  assign new_G5627 = ~new_G5621;
  assign new_G5630 = ~new_G5621 | ~new_G5628;
  assign new_G5715 = ~new_G5709;
  assign new_G5718 = ~new_G5709 | ~new_G5716;
  assign new_G6093 = ~new_G6087;
  assign new_G6096 = ~new_G6087 | ~new_G6094;
  assign new_G6151 = ~new_G6145;
  assign new_G6154 = ~new_G6145 | ~new_G6152;
  assign new_G6209 = ~new_G6203;
  assign new_G6212 = ~new_G6203 | ~new_G6210;
  assign new_G6301 = ~new_G6299 | ~new_G6300;
  assign new_G6961 = ~new_G6955;
  assign new_G6964 = ~new_G6955 | ~new_G6962;
  assign new_G7019 = ~new_G7013;
  assign new_G7022 = ~new_G7013 | ~new_G7020;
  assign new_G7081 = ~new_G7079 | ~new_G7080;
  assign new_G7169 = ~new_G7167 | ~new_G7168;
  assign G347 = new_G345 | new_G346;
  assign G350 = new_G348 | new_G349;
  assign G353 = new_G351 | new_G352;
  assign G356 = new_G354 | new_G355;
  assign new_G5059 = ~new_G5054 | ~new_G5057;
  assign new_G5147 = ~new_G5142 | ~new_G5145;
  assign new_G5629 = ~new_G5624 | ~new_G5627;
  assign new_G5717 = ~new_G5712 | ~new_G5715;
  assign new_G6095 = ~new_G6090 | ~new_G6093;
  assign new_G6153 = ~new_G6148 | ~new_G6151;
  assign new_G6211 = ~new_G6206 | ~new_G6209;
  assign new_G6963 = ~new_G6958 | ~new_G6961;
  assign new_G7021 = ~new_G7016 | ~new_G7019;
  assign new_G5061 = ~new_G5059 | ~new_G5060;
  assign new_G5149 = ~new_G5147 | ~new_G5148;
  assign new_G5511 = ~new_G5505;
  assign new_G5514 = ~new_G5505 | ~new_G5512;
  assign new_G5569 = ~new_G5563;
  assign new_G5572 = ~new_G5563 | ~new_G5570;
  assign new_G5631 = ~new_G5629 | ~new_G5630;
  assign new_G5719 = ~new_G5717 | ~new_G5718;
  assign new_G6097 = ~new_G6095 | ~new_G6096;
  assign new_G6155 = ~new_G6153 | ~new_G6154;
  assign new_G6213 = ~new_G6211 | ~new_G6212;
  assign new_G6307 = ~new_G6301;
  assign new_G6310 = ~new_G6301 | ~new_G6308;
  assign new_G6965 = ~new_G6963 | ~new_G6964;
  assign new_G7023 = ~new_G7021 | ~new_G7022;
  assign new_G7087 = ~new_G7081;
  assign new_G7090 = ~new_G7081 | ~new_G7088;
  assign new_G7175 = ~new_G7169;
  assign new_G7178 = ~new_G7169 | ~new_G7176;
  assign new_G5513 = ~new_G5508 | ~new_G5511;
  assign new_G5571 = ~new_G5566 | ~new_G5569;
  assign new_G6309 = ~new_G6304 | ~new_G6307;
  assign new_G7089 = ~new_G7084 | ~new_G7087;
  assign new_G7177 = ~new_G7172 | ~new_G7175;
  assign new_G5067 = ~new_G5061;
  assign new_G5070 = ~new_G5061 | ~new_G5068;
  assign new_G5155 = ~new_G5149;
  assign new_G5158 = ~new_G5149 | ~new_G5156;
  assign new_G5515 = ~new_G5513 | ~new_G5514;
  assign new_G5573 = ~new_G5571 | ~new_G5572;
  assign new_G5637 = ~new_G5631;
  assign new_G5640 = ~new_G5631 | ~new_G5638;
  assign new_G5725 = ~new_G5719;
  assign new_G5728 = ~new_G5719 | ~new_G5726;
  assign new_G6103 = ~new_G6097;
  assign new_G6106 = ~new_G6097 | ~new_G6104;
  assign new_G6161 = ~new_G6155;
  assign new_G6164 = ~new_G6155 | ~new_G6162;
  assign new_G6219 = ~new_G6213;
  assign new_G6222 = ~new_G6213 | ~new_G6220;
  assign new_G6311 = ~new_G6309 | ~new_G6310;
  assign new_G6971 = ~new_G6965;
  assign new_G6974 = ~new_G6965 | ~new_G6972;
  assign new_G7029 = ~new_G7023;
  assign new_G7032 = ~new_G7023 | ~new_G7030;
  assign new_G7091 = ~new_G7089 | ~new_G7090;
  assign new_G7179 = ~new_G7177 | ~new_G7178;
  assign new_G5069 = ~new_G5064 | ~new_G5067;
  assign new_G5157 = ~new_G5152 | ~new_G5155;
  assign new_G5639 = ~new_G5634 | ~new_G5637;
  assign new_G5727 = ~new_G5722 | ~new_G5725;
  assign new_G6105 = ~new_G6100 | ~new_G6103;
  assign new_G6163 = ~new_G6158 | ~new_G6161;
  assign new_G6221 = ~new_G6216 | ~new_G6219;
  assign new_G6973 = ~new_G6968 | ~new_G6971;
  assign new_G7031 = ~new_G7026 | ~new_G7029;
  assign new_G5521 = ~new_G5515;
  assign new_G1756 = ~new_G5515 | ~new_G5522;
  assign new_G5579 = ~new_G5573;
  assign new_G1761 = ~new_G5573 | ~new_G5580;
  assign new_G5071 = ~new_G5069 | ~new_G5070;
  assign new_G5159 = ~new_G5157 | ~new_G5158;
  assign new_G5641 = ~new_G5639 | ~new_G5640;
  assign new_G5729 = ~new_G5727 | ~new_G5728;
  assign new_G6107 = ~new_G6105 | ~new_G6106;
  assign new_G6165 = ~new_G6163 | ~new_G6164;
  assign new_G6223 = ~new_G6221 | ~new_G6222;
  assign new_G6317 = ~new_G6311;
  assign new_G6320 = ~new_G6311 | ~new_G6318;
  assign new_G6975 = ~new_G6973 | ~new_G6974;
  assign new_G7033 = ~new_G7031 | ~new_G7032;
  assign new_G7097 = ~new_G7091;
  assign new_G7100 = ~new_G7091 | ~new_G7098;
  assign new_G7185 = ~new_G7179;
  assign new_G7188 = ~new_G7179 | ~new_G7186;
  assign new_G1755 = ~new_G5518 | ~new_G5521;
  assign new_G1760 = ~new_G5576 | ~new_G5579;
  assign new_G6319 = ~new_G6314 | ~new_G6317;
  assign new_G7099 = ~new_G7094 | ~new_G7097;
  assign new_G7187 = ~new_G7182 | ~new_G7185;
  assign new_G1757 = ~new_G1755 | ~new_G1756;
  assign new_G1762 = ~new_G1760 | ~new_G1761;
  assign new_G6113 = ~new_G6107;
  assign new_G2818 = ~new_G6107 | ~new_G6114;
  assign new_G6171 = ~new_G6165;
  assign new_G2823 = ~new_G6165 | ~new_G6172;
  assign new_G6981 = ~new_G6975;
  assign new_G4058 = ~new_G6975 | ~new_G6982;
  assign new_G7039 = ~new_G7033;
  assign new_G4063 = ~new_G7033 | ~new_G7040;
  assign new_G5077 = ~new_G5071;
  assign new_G5080 = ~new_G5071 | ~new_G5078;
  assign new_G5165 = ~new_G5159;
  assign new_G5090 = ~new_G5159 | ~new_G5166;
  assign new_G5647 = ~new_G5641;
  assign new_G5650 = ~new_G5641 | ~new_G5648;
  assign new_G5735 = ~new_G5729;
  assign new_G5660 = ~new_G5729 | ~new_G5736;
  assign new_G6229 = ~new_G6223;
  assign new_G6232 = ~new_G6223 | ~new_G6230;
  assign new_G6321 = ~new_G6319 | ~new_G6320;
  assign new_G7101 = ~new_G7099 | ~new_G7100;
  assign new_G7189 = ~new_G7187 | ~new_G7188;
  assign new_G2817 = ~new_G6110 | ~new_G6113;
  assign new_G2822 = ~new_G6168 | ~new_G6171;
  assign new_G4057 = ~new_G6978 | ~new_G6981;
  assign new_G4062 = ~new_G7036 | ~new_G7039;
  assign new_G5079 = ~new_G5074 | ~new_G5077;
  assign new_G5089 = ~new_G5162 | ~new_G5165;
  assign new_G5649 = ~new_G5644 | ~new_G5647;
  assign new_G5659 = ~new_G5732 | ~new_G5735;
  assign new_G6231 = ~new_G6226 | ~new_G6229;
  assign new_G1782 = new_G1771 & new_G1762 & new_G1730;
  assign new_G1783 = new_G1771 & new_G1757 & new_G1726;
  assign new_G1784 = new_G1766 & new_G1762 & new_G1751;
  assign new_G1785 = new_G1766 & new_G1757 & new_G1754;
  assign new_G2819 = ~new_G2817 | ~new_G2818;
  assign new_G2824 = ~new_G2822 | ~new_G2823;
  assign new_G4059 = ~new_G4057 | ~new_G4058;
  assign new_G4064 = ~new_G4062 | ~new_G4063;
  assign new_G5081 = ~new_G5079 | ~new_G5080;
  assign new_G5091 = ~new_G5089 | ~new_G5090;
  assign new_G5651 = ~new_G5649 | ~new_G5650;
  assign new_G5661 = ~new_G5659 | ~new_G5660;
  assign new_G6233 = ~new_G6231 | ~new_G6232;
  assign new_G6327 = ~new_G6321;
  assign new_G6252 = ~new_G6321 | ~new_G6328;
  assign new_G7107 = ~new_G7101;
  assign new_G7110 = ~new_G7101 | ~new_G7108;
  assign new_G7195 = ~new_G7189;
  assign new_G7120 = ~new_G7189 | ~new_G7196;
  assign new_G5737 = new_G1785 | new_G1784 | new_G1782 | new_G1783;
  assign new_G6251 = ~new_G6324 | ~new_G6327;
  assign new_G7109 = ~new_G7104 | ~new_G7107;
  assign new_G7119 = ~new_G7192 | ~new_G7195;
  assign new_G5087 = ~new_G5081;
  assign new_G985 = ~new_G5081 | ~new_G5088;
  assign new_G5097 = ~new_G5091;
  assign new_G988 = ~new_G5091 | ~new_G5098;
  assign new_G5657 = ~new_G5651;
  assign new_G1776 = ~new_G5651 | ~new_G5658;
  assign new_G5667 = ~new_G5661;
  assign new_G1779 = ~new_G5661 | ~new_G5668;
  assign new_G2844 = new_G2833 & new_G2824 & new_G2784;
  assign new_G2845 = new_G2833 & new_G2819 & new_G2780;
  assign new_G2846 = new_G2828 & new_G2824 & new_G2813;
  assign new_G2847 = new_G2828 & new_G2819 & new_G2816;
  assign new_G4083 = new_G4072 & new_G4064 & new_G4032;
  assign new_G4084 = new_G4072 & new_G4059 & new_G4028;
  assign new_G4085 = new_G4067 & new_G4064 & new_G4053;
  assign new_G4086 = new_G4067 & new_G4059 & new_G4056;
  assign new_G6239 = ~new_G6233;
  assign new_G6242 = ~new_G6233 | ~new_G6240;
  assign new_G6253 = ~new_G6251 | ~new_G6252;
  assign new_G7111 = ~new_G7109 | ~new_G7110;
  assign new_G7121 = ~new_G7119 | ~new_G7120;
  assign new_G984 = ~new_G5084 | ~new_G5087;
  assign new_G987 = ~new_G5094 | ~new_G5097;
  assign new_G1775 = ~new_G5654 | ~new_G5657;
  assign new_G1778 = ~new_G5664 | ~new_G5667;
  assign new_G5743 = ~new_G5737;
  assign new_G6241 = ~new_G6236 | ~new_G6239;
  assign new_G6329 = new_G2847 | new_G2846 | new_G2844 | new_G2845;
  assign new_G7197 = new_G4086 | new_G4085 | new_G4083 | new_G4084;
  assign new_G986 = ~new_G984 | ~new_G985;
  assign new_G989 = ~new_G987 | ~new_G988;
  assign new_G1777 = ~new_G1775 | ~new_G1776;
  assign new_G1780 = ~new_G1778 | ~new_G1779;
  assign new_G6259 = ~new_G6253;
  assign new_G2841 = ~new_G6253 | ~new_G6260;
  assign new_G7117 = ~new_G7111;
  assign new_G4077 = ~new_G7111 | ~new_G7118;
  assign new_G7127 = ~new_G7121;
  assign new_G4080 = ~new_G7121 | ~new_G7128;
  assign new_G6243 = ~new_G6241 | ~new_G6242;
  assign new_G990 = ~new_G989;
  assign new_G996 = new_G975 & new_G986;
  assign new_G1781 = ~new_G1780;
  assign new_G1787 = new_G1766 & new_G1777;
  assign new_G2840 = ~new_G6256 | ~new_G6259;
  assign new_G6335 = ~new_G6329;
  assign new_G4076 = ~new_G7114 | ~new_G7117;
  assign new_G4079 = ~new_G7124 | ~new_G7127;
  assign new_G7203 = ~new_G7197;
  assign new_G995 = new_G990 & new_G980;
  assign new_G1786 = new_G1781 & new_G1771;
  assign new_G6249 = ~new_G6243;
  assign new_G2838 = ~new_G6243 | ~new_G6250;
  assign new_G2842 = ~new_G2840 | ~new_G2841;
  assign new_G4078 = ~new_G4076 | ~new_G4077;
  assign new_G4081 = ~new_G4079 | ~new_G4080;
  assign new_G2837 = ~new_G6246 | ~new_G6249;
  assign new_G2843 = ~new_G2842;
  assign new_G4082 = ~new_G4081;
  assign new_G4088 = new_G4067 & new_G4078;
  assign new_G5170 = new_G995 | new_G996;
  assign new_G5740 = new_G1786 | new_G1787;
  assign new_G2839 = ~new_G2837 | ~new_G2838;
  assign new_G2848 = new_G2843 & new_G2833;
  assign new_G4087 = new_G4082 & new_G4072;
  assign new_G1791 = ~new_G5740 | ~new_G5743;
  assign new_G1003 = ~new_G5170 | ~new_G5173;
  assign new_G5174 = ~new_G5170;
  assign new_G5744 = ~new_G5740;
  assign new_G2849 = new_G2828 & new_G2839;
  assign new_G7200 = new_G4087 | new_G4088;
  assign new_G1792 = ~new_G5737 | ~new_G5744;
  assign new_G1004 = ~new_G5167 | ~new_G5174;
  assign new_G6332 = new_G2848 | new_G2849;
  assign new_G320 = ~new_G1791 | ~new_G1792;
  assign new_G337 = ~new_G1003 | ~new_G1004;
  assign new_G4092 = ~new_G7200 | ~new_G7203;
  assign new_G7204 = ~new_G7200;
  assign G321 = ~new_G320;
  assign G338 = ~new_G337;
  assign new_G4093 = ~new_G7197 | ~new_G7204;
  assign new_G2855 = ~new_G6332 | ~new_G6335;
  assign new_G6336 = ~new_G6332;
  assign new_G369 = ~new_G4092 | ~new_G4093;
  assign new_G2856 = ~new_G6329 | ~new_G6336;
  assign G370 = ~new_G369;
  assign new_G398 = ~new_G2855 | ~new_G2856;
  assign G399 = ~new_G398;
endmodule
