// Benchmark "./benchmarks/iscas85/c1908" written by ABC on Sun Apr 28 12:32:37 2024

module c1908  ( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_G149, new_G153, new_G156, new_G160, new_G165, new_G168, new_G171,
    new_G175, new_G179, new_G184, new_G188, new_G191, new_G194, new_G198,
    new_G202, new_G206, new_G231, new_G233, new_G241, new_G244, new_G245,
    new_G248, new_G517, new_G529, new_G541, new_G553, new_G859, new_G862,
    new_G907, new_G909, new_G911, new_G918, new_G919, new_G922, new_G926,
    new_G930, new_G932, new_G934, new_G938, new_G943, new_G947, new_G949,
    new_G1506, new_G1514, new_G1522, new_G1530, new_G1538, new_G1546,
    new_G1554, new_G1562, new_G1570, new_G1578, new_G1586, new_G1594,
    new_G1602, new_G1610, new_G1618, new_G1626, new_G1512, new_G1520,
    new_G1528, new_G1536, new_G1544, new_G1552, new_G1560, new_G1568,
    new_G1576, new_G1584, new_G1592, new_G1600, new_G1608, new_G1616,
    new_G1624, new_G1632, new_G50, new_G52, new_G56, new_G58, new_G62,
    new_G64, new_G251, new_G254, new_G288, new_G291, new_G299, new_G302,
    new_G318, new_G321, new_G327, new_G330, new_G352, new_G355, new_G369,
    new_G382, new_G385, new_G853, new_G856, new_G893, new_G954, new_G955,
    new_G1050, new_G1053, new_G1176, new_G1179, new_G1197, new_G1207,
    new_G1222, new_G1244, new_G1278, new_G1290, new_G1300, new_G1312,
    new_G1332, new_G1335, new_G1442, new_G1450, new_G1458, new_G1466,
    new_G1474, new_G1482, new_G1490, new_G1498, new_G1634, new_G1644,
    new_G1657, new_G1665, new_G1697, new_G1705, new_G1713, new_G1721,
    new_G1745, new_G1753, new_G1785, new_G1793, new_G1814, new_G1817,
    new_G1830, new_G1833, new_G1841, new_G1849, new_G1854, new_G1857,
    new_G1870, new_G1873, new_G1878, new_G1881, new_G1642, new_G1652,
    new_G1056, new_G1057, new_G1182, new_G1183, new_G1211, new_G1298,
    new_G1320, new_G1338, new_G1339, new_G457, new_G459, new_G482,
    new_G487, new_G492, new_G505, new_G1456, new_G1448, new_G1472,
    new_G1464, new_G1488, new_G1480, new_G1504, new_G1496, new_G956,
    new_G967, new_G978, new_G979, new_G980, new_G1661, new_G990, new_G1669,
    new_G1030, new_G1701, new_G1040, new_G1709, new_G1058, new_G1717,
    new_G1068, new_G1725, new_G1078, new_G1090, new_G1100, new_G1749,
    new_G1112, new_G1757, new_G1154, new_G1789, new_G1166, new_G1797,
    new_G1194, new_G1201, new_G1204, new_G1820, new_G1821, new_G1230,
    new_G1836, new_G1837, new_G1252, new_G1256, new_G1845, new_G1268,
    new_G1853, new_G1860, new_G1861, new_G1286, new_G1876, new_G1877,
    new_G1308, new_G1884, new_G1885, new_G1654, new_G1662, new_G1694,
    new_G1702, new_G1710, new_G1718, new_G1726, new_G1734, new_G1742,
    new_G1750, new_G1782, new_G1790, new_G1838, new_G1846, new_G297,
    new_G298, new_G361, new_G362, new_G404, new_G405, new_G1225, new_G1226,
    new_G1247, new_G1248, new_G1281, new_G1282, new_G1303, new_G1304,
    new_G1315, new_G1316, new_G998, new_G988, new_G268, new_G1038,
    new_G1048, new_G1076, new_G1066, new_G1098, new_G1120, new_G1174,
    new_G363, new_G1210, new_G373, new_G1276, new_G406, new_G565, new_G566,
    new_G614, new_G615, new_G958, new_G969, new_G1660, new_G984, new_G1668,
    new_G994, new_G1700, new_G1034, new_G1708, new_G1044, new_G1716,
    new_G1062, new_G1724, new_G1072, new_G1732, new_G1086, new_G1740,
    new_G1748, new_G1104, new_G1108, new_G1756, new_G1116, new_G1788,
    new_G1158, new_G1162, new_G1796, new_G1170, new_G1200, new_G1203,
    new_G1227, new_G1249, new_G1844, new_G1260, new_G1264, new_G1852,
    new_G1272, new_G1283, new_G1305, new_G1317, new_G1410, new_G1418,
    new_G1426, new_G1434, new_G269, new_G372, new_G983, new_G993,
    new_G1033, new_G1043, new_G1061, new_G1071, new_G1103, new_G1115,
    new_G1157, new_G1169, new_G1184, new_G1202, new_G1259, new_G1271,
    new_G1322, new_G374, new_G396, new_G1321, new_G1424, new_G1416,
    new_G1440, new_G1432, new_G985, new_G995, new_G1035, new_G1045,
    new_G1063, new_G1073, new_G1105, new_G1117, new_G1159, new_G1171,
    new_G1212, new_G1231, new_G1232, new_G1253, new_G1254, new_G1261,
    new_G1273, new_G1287, new_G1288, new_G1309, new_G1310, new_G1192,
    new_G397, new_G1330, new_G1000, new_G1010, new_G1233, new_G1255,
    new_G1289, new_G1311, new_G1381, new_G257, new_G999, new_G260,
    new_G989, new_G272, new_G1039, new_G294, new_G1049, new_G305,
    new_G1077, new_G308, new_G1067, new_G333, new_G1121, new_G358,
    new_G1175, new_G1220, new_G388, new_G1277, new_G398, new_G1109,
    new_G1110, new_G1163, new_G1164, new_G1234, new_G1265, new_G1266,
    new_G1822, new_G1862, new_G1865, new_G258, new_G261, new_G273,
    new_G1018, new_G1008, new_G295, new_G306, new_G309, new_G334, new_G359,
    new_G389, new_G1385, new_G1111, new_G1165, new_G1267, new_G1886,
    new_G259, new_G262, new_G274, new_G296, new_G307, new_G310, new_G335,
    new_G360, new_G1242, new_G390, new_G1828, new_G1868, new_G1869,
    new_G1373, new_G1798, new_G1825, new_G265, new_G314, new_G336,
    new_G407, new_G1293, new_G1294, new_G1892, new_G1777, new_G1889,
    new_G410, new_G1377, new_G1804, new_G1237, new_G1829, new_G1295,
    new_G1670, new_G1678, new_G1729, new_G1737, new_G1761, new_G1769,
    new_G340, new_G343, new_G1781, new_G1238, new_G1325, new_G1893,
    new_G1340, new_G1352, new_G1673, new_G1681, new_G1801, new_G1897,
    new_G1905, new_G391, new_G1299, new_G1676, new_G1684, new_G1081,
    new_G1733, new_G1093, new_G1741, new_G1765, new_G1773, new_G1239,
    new_G1326, new_G1894, new_G1902, new_G392, new_G1360, new_G1003,
    new_G1677, new_G1013, new_G1685, new_G1082, new_G1094, new_G1122,
    new_G1134, new_G1187, new_G1805, new_G1327, new_G1901, new_G1348,
    new_G1909, new_G1758, new_G1766, new_G377, new_G1243, new_G393,
    new_G1004, new_G1014, new_G1083, new_G1095, new_G1188, new_G1900,
    new_G1344, new_G1908, new_G1356, new_G1142, new_G378, new_G399,
    new_G1331, new_G1005, new_G1015, new_G1764, new_G1126, new_G1130,
    new_G1772, new_G1138, new_G1189, new_G1343, new_G1355, new_G324,
    new_G1099, new_G379, new_G400, new_G449, new_G1087, new_G1088,
    new_G1125, new_G1137, new_G1345, new_G1357, new_G1397, new_G277,
    new_G1019, new_G280, new_G1009, new_G325, new_G364, new_G1193,
    new_G401, new_G1089, new_G1127, new_G1139, new_G278, new_G281,
    new_G326, new_G365, new_G413, new_G1361, new_G1401, new_G445,
    new_G1349, new_G1350, new_G1389, new_G1493, new_G1501, new_G1689,
    new_G279, new_G282, new_G346, new_G1143, new_G366, new_G414, new_G453,
    new_G1131, new_G1132, new_G1351, new_G1365, new_G1405, new_G285,
    new_G347, new_G367, new_G415, new_G1393, new_G556, new_G1505, new_G559,
    new_G1497, new_G1693, new_G1133, new_G1477, new_G1485, new_G1809,
    new_G348, new_G1369, new_G1409, new_G557, new_G560, new_G1362,
    new_G1378, new_G1429, new_G1437, new_G1686, new_G1774, new_G1910,
    new_G1918, new_G544, new_G1489, new_G547, new_G1481, new_G558,
    new_G561, new_G1813, new_G1370, new_G1368, new_G417, new_G1384,
    new_G424, new_G508, new_G1441, new_G511, new_G1433, new_G545, new_G548,
    new_G564, new_G1692, new_G1024, new_G1780, new_G1148, new_G1916,
    new_G1924, new_G416, new_G1376, new_G421, new_G423, new_G509, new_G512,
    new_G546, new_G549, new_G719, new_G722, new_G1023, new_G1147, new_G418,
    new_G420, new_G425, new_G510, new_G513, new_G552, new_G1025, new_G1149,
    new_G419, new_G422, new_G441, new_G516, new_G725, new_G728, new_G1029,
    new_G1153, new_G433, new_G437, new_G663, new_G666, new_G731, new_G746,
    new_G756, new_G770, new_G1461, new_G1469, new_G1413, new_G1421,
    new_G1445, new_G1453, new_G532, new_G1473, new_G535, new_G1465,
    new_G495, new_G1425, new_G498, new_G1417, new_G520, new_G1457,
    new_G523, new_G1449, new_G533, new_G536, new_G496, new_G499, new_G521,
    new_G524, new_G534, new_G537, new_G497, new_G500, new_G522, new_G525,
    new_G540, new_G503, new_G528, new_G669, new_G672, new_G569, new_G588,
    new_G618, new_G639, new_G867, new_G588a, new_G588b, new_G639a,
    new_G639b, new_G675, new_G688, new_G696, new_G710, new_G73, new_G572,
    new_G573, new_G621, new_G622, new_G776, new_G780, new_G784, new_G788,
    new_G812, new_G832, new_G836, new_G1509, new_G1517, new_G1525,
    new_G1533, new_G1581, new_G1621, new_G1629, new_G792, new_G796,
    new_G800, new_G804, new_G808, new_G816, new_G820, new_G824, new_G828,
    new_G871, new_G873, new_G875, new_G877, new_G879, new_G881, new_G883,
    new_G885, new_G1541, new_G1549, new_G1557, new_G1565, new_G1573,
    new_G1589, new_G1597, new_G1605, new_G1613, new_G1, new_G1513, new_G4,
    new_G1521, new_G7, new_G1529, new_G10, new_G1537, new_G28, new_G1585,
    new_G43, new_G1625, new_G46, new_G1633, new_G886, new_G2, new_G5,
    new_G8, new_G11, new_G13, new_G1545, new_G16, new_G1553, new_G19,
    new_G1561, new_G22, new_G1569, new_G25, new_G1577, new_G29, new_G31,
    new_G1593, new_G34, new_G1601, new_G37, new_G1609, new_G40, new_G1617,
    new_G44, new_G47, new_G857, new_G860, new_G863, new_G865, new_G14,
    new_G17, new_G20, new_G23, new_G26, new_G32, new_G35, new_G38, new_G41,
    new_G1913, new_G1921, new_G887, new_G462, new_G74, new_G1637,
    new_G1917, new_G1647, new_G1925, new_G1020, new_G1144, new_G1386,
    new_G1394, new_G1402, new_G1638, new_G1648, new_G1806, new_G1639,
    new_G1649, new_G287, new_G350, new_G427, new_G429, new_G431, new_G1028,
    new_G1152, new_G1392, new_G1400, new_G1408, new_G1812, new_G1216,
    new_G286, new_G349, new_G426, new_G428, new_G430, new_G67, new_G1643,
    new_G70, new_G1653, new_G1215, new_G49, new_G53, new_G59, new_G61,
    new_G65, new_G68, new_G71, new_G1217, new_G375, new_G1221, new_G376,
    new_G55;
  assign new_G149 = ~G101;
  assign new_G153 = ~G104;
  assign new_G156 = ~G107;
  assign new_G160 = ~G110;
  assign new_G165 = ~G113;
  assign new_G168 = ~G116;
  assign new_G171 = ~G119;
  assign new_G175 = ~G122;
  assign new_G179 = ~G125;
  assign new_G184 = ~G128;
  assign new_G188 = ~G131;
  assign new_G191 = ~G134;
  assign new_G194 = ~G137;
  assign new_G198 = ~G140;
  assign new_G202 = ~G143;
  assign new_G206 = ~G146;
  assign new_G231 = ~G224 | ~G898;
  assign new_G233 = ~G227 | ~G900;
  assign new_G241 = ~G237;
  assign new_G244 = ~G237;
  assign new_G245 = G234;
  assign new_G248 = G234;
  assign new_G517 = ~G469;
  assign new_G529 = ~G472;
  assign new_G541 = ~G475;
  assign new_G553 = ~G478;
  assign new_G859 = ~G953;
  assign new_G862 = ~G953;
  assign new_G907 = ~G898;
  assign new_G909 = ~G900;
  assign new_G911 = G902;
  assign new_G918 = ~G902;
  assign new_G919 = G902;
  assign new_G922 = ~G902;
  assign new_G926 = G952;
  assign new_G930 = ~G952;
  assign new_G932 = ~G952;
  assign new_G934 = G953;
  assign new_G938 = ~G953;
  assign new_G943 = G953;
  assign new_G947 = G953;
  assign new_G949 = ~G953;
  assign new_G1506 = G101;
  assign new_G1514 = G104;
  assign new_G1522 = G107;
  assign new_G1530 = G110;
  assign new_G1538 = G113;
  assign new_G1546 = G116;
  assign new_G1554 = G119;
  assign new_G1562 = G122;
  assign new_G1570 = G125;
  assign new_G1578 = G128;
  assign new_G1586 = G131;
  assign new_G1594 = G134;
  assign new_G1602 = G137;
  assign new_G1610 = G140;
  assign new_G1618 = G143;
  assign new_G1626 = G146;
  assign new_G1512 = ~new_G1506;
  assign new_G1520 = ~new_G1514;
  assign new_G1528 = ~new_G1522;
  assign new_G1536 = ~new_G1530;
  assign new_G1544 = ~new_G1538;
  assign new_G1552 = ~new_G1546;
  assign new_G1560 = ~new_G1554;
  assign new_G1568 = ~new_G1562;
  assign new_G1576 = ~new_G1570;
  assign new_G1584 = ~new_G1578;
  assign new_G1592 = ~new_G1586;
  assign new_G1600 = ~new_G1594;
  assign new_G1608 = ~new_G1602;
  assign new_G1616 = ~new_G1610;
  assign new_G1624 = ~new_G1618;
  assign new_G1632 = ~new_G1626;
  assign new_G50 = ~new_G930 | ~new_G947;
  assign new_G52 = ~new_G930 | ~new_G947;
  assign new_G56 = ~new_G930 | ~new_G947;
  assign new_G58 = ~new_G930 | ~new_G947;
  assign new_G62 = ~new_G930 | ~new_G947;
  assign new_G64 = ~new_G930 | ~new_G947;
  assign new_G251 = new_G149;
  assign new_G254 = new_G153;
  assign new_G288 = new_G165;
  assign new_G291 = new_G168;
  assign new_G299 = new_G184;
  assign new_G302 = new_G202;
  assign new_G318 = G224 & new_G938;
  assign new_G321 = new_G179;
  assign new_G327 = new_G188;
  assign new_G330 = new_G191;
  assign new_G352 = G227 & new_G938;
  assign new_G355 = new_G198;
  assign new_G369 = new_G938 & G210 & new_G241;
  assign new_G382 = new_G206;
  assign new_G385 = new_G198;
  assign new_G853 = ~new_G943 | ~new_G907;
  assign new_G856 = ~new_G943 | ~new_G909;
  assign new_G893 = ~new_G248 | ~G237;
  assign new_G954 = ~new_G248 | ~new_G922;
  assign new_G955 = ~new_G244 | ~new_G922;
  assign new_G1050 = new_G160;
  assign new_G1053 = new_G175;
  assign new_G1176 = new_G179;
  assign new_G1179 = new_G198;
  assign new_G1197 = new_G149;
  assign new_G1207 = new_G149;
  assign new_G1222 = new_G153;
  assign new_G1244 = new_G188;
  assign new_G1278 = new_G156;
  assign new_G1290 = new_G938 & G217 & new_G245;
  assign new_G1300 = new_G191;
  assign new_G1312 = new_G160;
  assign new_G1332 = new_G194;
  assign new_G1335 = new_G938 & G221 & new_G245;
  assign new_G1442 = new_G517;
  assign new_G1450 = new_G517;
  assign new_G1458 = new_G529;
  assign new_G1466 = new_G529;
  assign new_G1474 = new_G541;
  assign new_G1482 = new_G541;
  assign new_G1490 = new_G553;
  assign new_G1498 = new_G553;
  assign new_G1634 = new_G231 & new_G934;
  assign new_G1644 = new_G233 & new_G934;
  assign new_G1657 = new_G156;
  assign new_G1665 = new_G156;
  assign new_G1697 = new_G171;
  assign new_G1705 = new_G171;
  assign new_G1713 = new_G206;
  assign new_G1721 = new_G206;
  assign new_G1745 = new_G194;
  assign new_G1753 = new_G194;
  assign new_G1785 = new_G160;
  assign new_G1793 = new_G160;
  assign new_G1814 = new_G165;
  assign new_G1817 = new_G175;
  assign new_G1830 = new_G938 & G214 & new_G241;
  assign new_G1833 = new_G202;
  assign new_G1841 = new_G179;
  assign new_G1849 = new_G179;
  assign new_G1854 = new_G168;
  assign new_G1857 = new_G175;
  assign new_G1870 = new_G184;
  assign new_G1873 = new_G202;
  assign new_G1878 = new_G171;
  assign new_G1881 = new_G184;
  assign new_G1642 = ~new_G1634;
  assign new_G1652 = ~new_G1644;
  assign new_G1056 = ~new_G1050;
  assign new_G1057 = ~new_G1053;
  assign new_G1182 = ~new_G1176;
  assign new_G1183 = ~new_G1179;
  assign new_G1211 = ~new_G1207;
  assign new_G1298 = ~new_G1290;
  assign new_G1320 = ~new_G1312;
  assign new_G1338 = ~new_G1332;
  assign new_G1339 = ~new_G1335;
  assign new_G457 = G210 & new_G955;
  assign new_G459 = G217 & new_G954;
  assign new_G482 = ~G214 | ~new_G955;
  assign new_G487 = ~G221 | ~new_G954;
  assign new_G492 = ~G210 | ~new_G955;
  assign new_G505 = ~G217 | ~new_G954;
  assign new_G1456 = ~new_G1450;
  assign new_G1448 = ~new_G1442;
  assign new_G1472 = ~new_G1466;
  assign new_G1464 = ~new_G1458;
  assign new_G1488 = ~new_G1482;
  assign new_G1480 = ~new_G1474;
  assign new_G1504 = ~new_G1498;
  assign new_G1496 = ~new_G1490;
  assign new_G956 = ~new_G893 | ~new_G943 | ~new_G907 | ~new_G919;
  assign new_G967 = ~new_G893 | ~new_G943 | ~new_G909 | ~new_G919;
  assign new_G978 = ~new_G893 | ~new_G926 | ~new_G949;
  assign new_G979 = new_G893 & new_G926 & new_G949;
  assign new_G980 = new_G251;
  assign new_G1661 = ~new_G1657;
  assign new_G990 = new_G251;
  assign new_G1669 = ~new_G1665;
  assign new_G1030 = new_G288;
  assign new_G1701 = ~new_G1697;
  assign new_G1040 = new_G288;
  assign new_G1709 = ~new_G1705;
  assign new_G1058 = new_G299;
  assign new_G1717 = ~new_G1713;
  assign new_G1068 = new_G299;
  assign new_G1725 = ~new_G1721;
  assign new_G1078 = new_G318;
  assign new_G1090 = new_G318;
  assign new_G1100 = new_G327;
  assign new_G1749 = ~new_G1745;
  assign new_G1112 = new_G327;
  assign new_G1757 = ~new_G1753;
  assign new_G1154 = new_G352;
  assign new_G1789 = ~new_G1785;
  assign new_G1166 = new_G352;
  assign new_G1797 = ~new_G1793;
  assign new_G1194 = new_G369;
  assign new_G1201 = ~new_G1197;
  assign new_G1204 = new_G369;
  assign new_G1820 = ~new_G1814;
  assign new_G1821 = ~new_G1817;
  assign new_G1230 = ~new_G1222;
  assign new_G1836 = ~new_G1830;
  assign new_G1837 = ~new_G1833;
  assign new_G1252 = ~new_G1244;
  assign new_G1256 = new_G382;
  assign new_G1845 = ~new_G1841;
  assign new_G1268 = new_G382;
  assign new_G1853 = ~new_G1849;
  assign new_G1860 = ~new_G1854;
  assign new_G1861 = ~new_G1857;
  assign new_G1286 = ~new_G1278;
  assign new_G1876 = ~new_G1870;
  assign new_G1877 = ~new_G1873;
  assign new_G1308 = ~new_G1300;
  assign new_G1884 = ~new_G1878;
  assign new_G1885 = ~new_G1881;
  assign new_G1654 = new_G254;
  assign new_G1662 = new_G254;
  assign new_G1694 = new_G291;
  assign new_G1702 = new_G291;
  assign new_G1710 = new_G302;
  assign new_G1718 = new_G302;
  assign new_G1726 = new_G321;
  assign new_G1734 = new_G321;
  assign new_G1742 = new_G330;
  assign new_G1750 = new_G330;
  assign new_G1782 = new_G355;
  assign new_G1790 = new_G355;
  assign new_G1838 = new_G385;
  assign new_G1846 = new_G385;
  assign new_G297 = ~new_G1053 | ~new_G1056;
  assign new_G298 = ~new_G1050 | ~new_G1057;
  assign new_G361 = ~new_G1179 | ~new_G1182;
  assign new_G362 = ~new_G1176 | ~new_G1183;
  assign new_G404 = ~new_G1335 | ~new_G1338;
  assign new_G405 = ~new_G1332 | ~new_G1339;
  assign new_G1225 = ~new_G1817 | ~new_G1820;
  assign new_G1226 = ~new_G1814 | ~new_G1821;
  assign new_G1247 = ~new_G1833 | ~new_G1836;
  assign new_G1248 = ~new_G1830 | ~new_G1837;
  assign new_G1281 = ~new_G1857 | ~new_G1860;
  assign new_G1282 = ~new_G1854 | ~new_G1861;
  assign new_G1303 = ~new_G1873 | ~new_G1876;
  assign new_G1304 = ~new_G1870 | ~new_G1877;
  assign new_G1315 = ~new_G1881 | ~new_G1884;
  assign new_G1316 = ~new_G1878 | ~new_G1885;
  assign new_G998 = ~new_G990;
  assign new_G988 = ~new_G980;
  assign new_G268 = ~new_G297 | ~new_G298;
  assign new_G1038 = ~new_G1030;
  assign new_G1048 = ~new_G1040;
  assign new_G1076 = ~new_G1068;
  assign new_G1066 = ~new_G1058;
  assign new_G1098 = ~new_G1090;
  assign new_G1120 = ~new_G1112;
  assign new_G1174 = ~new_G1166;
  assign new_G363 = ~new_G361 | ~new_G362;
  assign new_G1210 = ~new_G1204;
  assign new_G373 = ~new_G1204 | ~new_G1211;
  assign new_G1276 = ~new_G1268;
  assign new_G406 = ~new_G404 | ~new_G405;
  assign new_G565 = ~new_G482;
  assign new_G566 = new_G482;
  assign new_G614 = ~new_G487;
  assign new_G615 = new_G487;
  assign new_G958 = ~new_G956 | ~new_G978;
  assign new_G969 = ~new_G967 | ~new_G978;
  assign new_G1660 = ~new_G1654;
  assign new_G984 = ~new_G1654 | ~new_G1661;
  assign new_G1668 = ~new_G1662;
  assign new_G994 = ~new_G1662 | ~new_G1669;
  assign new_G1700 = ~new_G1694;
  assign new_G1034 = ~new_G1694 | ~new_G1701;
  assign new_G1708 = ~new_G1702;
  assign new_G1044 = ~new_G1702 | ~new_G1709;
  assign new_G1716 = ~new_G1710;
  assign new_G1062 = ~new_G1710 | ~new_G1717;
  assign new_G1724 = ~new_G1718;
  assign new_G1072 = ~new_G1718 | ~new_G1725;
  assign new_G1732 = ~new_G1726;
  assign new_G1086 = ~new_G1078;
  assign new_G1740 = ~new_G1734;
  assign new_G1748 = ~new_G1742;
  assign new_G1104 = ~new_G1742 | ~new_G1749;
  assign new_G1108 = ~new_G1100;
  assign new_G1756 = ~new_G1750;
  assign new_G1116 = ~new_G1750 | ~new_G1757;
  assign new_G1788 = ~new_G1782;
  assign new_G1158 = ~new_G1782 | ~new_G1789;
  assign new_G1162 = ~new_G1154;
  assign new_G1796 = ~new_G1790;
  assign new_G1170 = ~new_G1790 | ~new_G1797;
  assign new_G1200 = ~new_G1194;
  assign new_G1203 = ~new_G1194 | ~new_G1201;
  assign new_G1227 = ~new_G1225 | ~new_G1226;
  assign new_G1249 = ~new_G1247 | ~new_G1248;
  assign new_G1844 = ~new_G1838;
  assign new_G1260 = ~new_G1838 | ~new_G1845;
  assign new_G1264 = ~new_G1256;
  assign new_G1852 = ~new_G1846;
  assign new_G1272 = ~new_G1846 | ~new_G1853;
  assign new_G1283 = ~new_G1281 | ~new_G1282;
  assign new_G1305 = ~new_G1303 | ~new_G1304;
  assign new_G1317 = ~new_G1315 | ~new_G1316;
  assign new_G1410 = new_G492;
  assign new_G1418 = new_G492;
  assign new_G1426 = new_G505;
  assign new_G1434 = new_G505;
  assign new_G269 = ~new_G268;
  assign new_G372 = ~new_G1207 | ~new_G1210;
  assign new_G983 = ~new_G1657 | ~new_G1660;
  assign new_G993 = ~new_G1665 | ~new_G1668;
  assign new_G1033 = ~new_G1697 | ~new_G1700;
  assign new_G1043 = ~new_G1705 | ~new_G1708;
  assign new_G1061 = ~new_G1713 | ~new_G1716;
  assign new_G1071 = ~new_G1721 | ~new_G1724;
  assign new_G1103 = ~new_G1745 | ~new_G1748;
  assign new_G1115 = ~new_G1753 | ~new_G1756;
  assign new_G1157 = ~new_G1785 | ~new_G1788;
  assign new_G1169 = ~new_G1793 | ~new_G1796;
  assign new_G1184 = ~new_G363;
  assign new_G1202 = ~new_G1197 | ~new_G1200;
  assign new_G1259 = ~new_G1841 | ~new_G1844;
  assign new_G1271 = ~new_G1849 | ~new_G1852;
  assign new_G1322 = ~new_G406;
  assign new_G374 = ~new_G372 | ~new_G373;
  assign new_G396 = ~new_G1317 | ~new_G1320;
  assign new_G1321 = ~new_G1317;
  assign new_G1424 = ~new_G1418;
  assign new_G1416 = ~new_G1410;
  assign new_G1440 = ~new_G1434;
  assign new_G1432 = ~new_G1426;
  assign new_G985 = ~new_G983 | ~new_G984;
  assign new_G995 = ~new_G993 | ~new_G994;
  assign new_G1035 = ~new_G1033 | ~new_G1034;
  assign new_G1045 = ~new_G1043 | ~new_G1044;
  assign new_G1063 = ~new_G1061 | ~new_G1062;
  assign new_G1073 = ~new_G1071 | ~new_G1072;
  assign new_G1105 = ~new_G1103 | ~new_G1104;
  assign new_G1117 = ~new_G1115 | ~new_G1116;
  assign new_G1159 = ~new_G1157 | ~new_G1158;
  assign new_G1171 = ~new_G1169 | ~new_G1170;
  assign new_G1212 = ~new_G1202 | ~new_G1203;
  assign new_G1231 = ~new_G1227;
  assign new_G1232 = ~new_G1227 | ~new_G1230;
  assign new_G1253 = ~new_G1249;
  assign new_G1254 = ~new_G1249 | ~new_G1252;
  assign new_G1261 = ~new_G1259 | ~new_G1260;
  assign new_G1273 = ~new_G1271 | ~new_G1272;
  assign new_G1287 = ~new_G1283;
  assign new_G1288 = ~new_G1283 | ~new_G1286;
  assign new_G1309 = ~new_G1305;
  assign new_G1310 = ~new_G1305 | ~new_G1308;
  assign new_G1192 = ~new_G1184;
  assign new_G397 = ~new_G1312 | ~new_G1321;
  assign new_G1330 = ~new_G1322;
  assign new_G1000 = new_G269;
  assign new_G1010 = new_G269;
  assign new_G1233 = ~new_G1222 | ~new_G1231;
  assign new_G1255 = ~new_G1244 | ~new_G1253;
  assign new_G1289 = ~new_G1278 | ~new_G1287;
  assign new_G1311 = ~new_G1300 | ~new_G1309;
  assign new_G1381 = ~new_G374;
  assign new_G257 = ~new_G995 | ~new_G998;
  assign new_G999 = ~new_G995;
  assign new_G260 = ~new_G985 | ~new_G988;
  assign new_G989 = ~new_G985;
  assign new_G272 = ~new_G1035 | ~new_G1038;
  assign new_G1039 = ~new_G1035;
  assign new_G294 = ~new_G1045 | ~new_G1048;
  assign new_G1049 = ~new_G1045;
  assign new_G305 = ~new_G1073 | ~new_G1076;
  assign new_G1077 = ~new_G1073;
  assign new_G308 = ~new_G1063 | ~new_G1066;
  assign new_G1067 = ~new_G1063;
  assign new_G333 = ~new_G1117 | ~new_G1120;
  assign new_G1121 = ~new_G1117;
  assign new_G358 = ~new_G1171 | ~new_G1174;
  assign new_G1175 = ~new_G1171;
  assign new_G1220 = ~new_G1212;
  assign new_G388 = ~new_G1273 | ~new_G1276;
  assign new_G1277 = ~new_G1273;
  assign new_G398 = ~new_G396 | ~new_G397;
  assign new_G1109 = ~new_G1105;
  assign new_G1110 = ~new_G1105 | ~new_G1108;
  assign new_G1163 = ~new_G1159;
  assign new_G1164 = ~new_G1159 | ~new_G1162;
  assign new_G1234 = ~new_G1232 | ~new_G1233;
  assign new_G1265 = ~new_G1261;
  assign new_G1266 = ~new_G1261 | ~new_G1264;
  assign new_G1822 = ~new_G1254 | ~new_G1255;
  assign new_G1862 = ~new_G1310 | ~new_G1311;
  assign new_G1865 = ~new_G1288 | ~new_G1289;
  assign new_G258 = ~new_G990 | ~new_G999;
  assign new_G261 = ~new_G980 | ~new_G989;
  assign new_G273 = ~new_G1030 | ~new_G1039;
  assign new_G1018 = ~new_G1010;
  assign new_G1008 = ~new_G1000;
  assign new_G295 = ~new_G1040 | ~new_G1049;
  assign new_G306 = ~new_G1068 | ~new_G1077;
  assign new_G309 = ~new_G1058 | ~new_G1067;
  assign new_G334 = ~new_G1112 | ~new_G1121;
  assign new_G359 = ~new_G1166 | ~new_G1175;
  assign new_G389 = ~new_G1268 | ~new_G1277;
  assign new_G1385 = ~new_G1381;
  assign new_G1111 = ~new_G1100 | ~new_G1109;
  assign new_G1165 = ~new_G1154 | ~new_G1163;
  assign new_G1267 = ~new_G1256 | ~new_G1265;
  assign new_G1886 = ~new_G398;
  assign new_G259 = ~new_G257 | ~new_G258;
  assign new_G262 = ~new_G260 | ~new_G261;
  assign new_G274 = ~new_G272 | ~new_G273;
  assign new_G296 = ~new_G294 | ~new_G295;
  assign new_G307 = ~new_G305 | ~new_G306;
  assign new_G310 = ~new_G308 | ~new_G309;
  assign new_G335 = ~new_G333 | ~new_G334;
  assign new_G360 = ~new_G358 | ~new_G359;
  assign new_G1242 = ~new_G1234;
  assign new_G390 = ~new_G388 | ~new_G389;
  assign new_G1828 = ~new_G1822;
  assign new_G1868 = ~new_G1862;
  assign new_G1869 = ~new_G1865;
  assign new_G1373 = ~new_G1164 | ~new_G1165;
  assign new_G1798 = ~new_G1110 | ~new_G1111;
  assign new_G1825 = ~new_G1266 | ~new_G1267;
  assign new_G265 = ~new_G259;
  assign new_G314 = ~new_G307;
  assign new_G336 = ~new_G335;
  assign new_G407 = ~new_G296;
  assign new_G1293 = ~new_G1865 | ~new_G1868;
  assign new_G1294 = ~new_G1862 | ~new_G1869;
  assign new_G1892 = ~new_G1886;
  assign new_G1777 = ~new_G360;
  assign new_G1889 = ~new_G390;
  assign new_G410 = new_G310;
  assign new_G1377 = ~new_G1373;
  assign new_G1804 = ~new_G1798;
  assign new_G1237 = ~new_G1825 | ~new_G1828;
  assign new_G1829 = ~new_G1825;
  assign new_G1295 = ~new_G1293 | ~new_G1294;
  assign new_G1670 = new_G274;
  assign new_G1678 = new_G274;
  assign new_G1729 = new_G310;
  assign new_G1737 = new_G310;
  assign new_G1761 = new_G262;
  assign new_G1769 = new_G262;
  assign new_G340 = new_G336;
  assign new_G343 = new_G314;
  assign new_G1781 = ~new_G1777;
  assign new_G1238 = ~new_G1822 | ~new_G1829;
  assign new_G1325 = ~new_G1889 | ~new_G1892;
  assign new_G1893 = ~new_G1889;
  assign new_G1340 = new_G407;
  assign new_G1352 = new_G407;
  assign new_G1673 = new_G265;
  assign new_G1681 = new_G265;
  assign new_G1801 = new_G314;
  assign new_G1897 = new_G336;
  assign new_G1905 = new_G336;
  assign new_G391 = ~new_G1295 | ~new_G1298;
  assign new_G1299 = ~new_G1295;
  assign new_G1676 = ~new_G1670;
  assign new_G1684 = ~new_G1678;
  assign new_G1081 = ~new_G1729 | ~new_G1732;
  assign new_G1733 = ~new_G1729;
  assign new_G1093 = ~new_G1737 | ~new_G1740;
  assign new_G1741 = ~new_G1737;
  assign new_G1765 = ~new_G1761;
  assign new_G1773 = ~new_G1769;
  assign new_G1239 = ~new_G1237 | ~new_G1238;
  assign new_G1326 = ~new_G1886 | ~new_G1893;
  assign new_G1894 = new_G410;
  assign new_G1902 = new_G410;
  assign new_G392 = ~new_G1290 | ~new_G1299;
  assign new_G1360 = ~new_G1352;
  assign new_G1003 = ~new_G1673 | ~new_G1676;
  assign new_G1677 = ~new_G1673;
  assign new_G1013 = ~new_G1681 | ~new_G1684;
  assign new_G1685 = ~new_G1681;
  assign new_G1082 = ~new_G1726 | ~new_G1733;
  assign new_G1094 = ~new_G1734 | ~new_G1741;
  assign new_G1122 = new_G340;
  assign new_G1134 = new_G340;
  assign new_G1187 = ~new_G1801 | ~new_G1804;
  assign new_G1805 = ~new_G1801;
  assign new_G1327 = ~new_G1325 | ~new_G1326;
  assign new_G1901 = ~new_G1897;
  assign new_G1348 = ~new_G1340;
  assign new_G1909 = ~new_G1905;
  assign new_G1758 = new_G343;
  assign new_G1766 = new_G343;
  assign new_G377 = ~new_G1239 | ~new_G1242;
  assign new_G1243 = ~new_G1239;
  assign new_G393 = ~new_G391 | ~new_G392;
  assign new_G1004 = ~new_G1670 | ~new_G1677;
  assign new_G1014 = ~new_G1678 | ~new_G1685;
  assign new_G1083 = ~new_G1081 | ~new_G1082;
  assign new_G1095 = ~new_G1093 | ~new_G1094;
  assign new_G1188 = ~new_G1798 | ~new_G1805;
  assign new_G1900 = ~new_G1894;
  assign new_G1344 = ~new_G1894 | ~new_G1901;
  assign new_G1908 = ~new_G1902;
  assign new_G1356 = ~new_G1902 | ~new_G1909;
  assign new_G1142 = ~new_G1134;
  assign new_G378 = ~new_G1234 | ~new_G1243;
  assign new_G399 = ~new_G1327 | ~new_G1330;
  assign new_G1331 = ~new_G1327;
  assign new_G1005 = ~new_G1003 | ~new_G1004;
  assign new_G1015 = ~new_G1013 | ~new_G1014;
  assign new_G1764 = ~new_G1758;
  assign new_G1126 = ~new_G1758 | ~new_G1765;
  assign new_G1130 = ~new_G1122;
  assign new_G1772 = ~new_G1766;
  assign new_G1138 = ~new_G1766 | ~new_G1773;
  assign new_G1189 = ~new_G1187 | ~new_G1188;
  assign new_G1343 = ~new_G1897 | ~new_G1900;
  assign new_G1355 = ~new_G1905 | ~new_G1908;
  assign new_G324 = ~new_G1095 | ~new_G1098;
  assign new_G1099 = ~new_G1095;
  assign new_G379 = ~new_G377 | ~new_G378;
  assign new_G400 = ~new_G1322 | ~new_G1331;
  assign new_G449 = ~new_G393 | ~new_G918;
  assign new_G1087 = ~new_G1083;
  assign new_G1088 = ~new_G1083 | ~new_G1086;
  assign new_G1125 = ~new_G1761 | ~new_G1764;
  assign new_G1137 = ~new_G1769 | ~new_G1772;
  assign new_G1345 = ~new_G1343 | ~new_G1344;
  assign new_G1357 = ~new_G1355 | ~new_G1356;
  assign new_G1397 = new_G393;
  assign new_G277 = ~new_G1015 | ~new_G1018;
  assign new_G1019 = ~new_G1015;
  assign new_G280 = ~new_G1005 | ~new_G1008;
  assign new_G1009 = ~new_G1005;
  assign new_G325 = ~new_G1090 | ~new_G1099;
  assign new_G364 = ~new_G1189 | ~new_G1192;
  assign new_G1193 = ~new_G1189;
  assign new_G401 = ~new_G399 | ~new_G400;
  assign new_G1089 = ~new_G1078 | ~new_G1087;
  assign new_G1127 = ~new_G1125 | ~new_G1126;
  assign new_G1139 = ~new_G1137 | ~new_G1138;
  assign new_G278 = ~new_G1010 | ~new_G1019;
  assign new_G281 = ~new_G1000 | ~new_G1009;
  assign new_G326 = ~new_G324 | ~new_G325;
  assign new_G365 = ~new_G1184 | ~new_G1193;
  assign new_G413 = ~new_G1357 | ~new_G1360;
  assign new_G1361 = ~new_G1357;
  assign new_G1401 = ~new_G1397;
  assign new_G445 = ~new_G379 | ~new_G918;
  assign new_G1349 = ~new_G1345;
  assign new_G1350 = ~new_G1345 | ~new_G1348;
  assign new_G1389 = new_G379;
  assign new_G1493 = new_G449;
  assign new_G1501 = new_G449;
  assign new_G1689 = ~new_G1088 | ~new_G1089;
  assign new_G279 = ~new_G277 | ~new_G278;
  assign new_G282 = ~new_G280 | ~new_G281;
  assign new_G346 = ~new_G1139 | ~new_G1142;
  assign new_G1143 = ~new_G1139;
  assign new_G366 = ~new_G364 | ~new_G365;
  assign new_G414 = ~new_G1352 | ~new_G1361;
  assign new_G453 = ~new_G401 | ~new_G918;
  assign new_G1131 = ~new_G1127;
  assign new_G1132 = ~new_G1127 | ~new_G1130;
  assign new_G1351 = ~new_G1340 | ~new_G1349;
  assign new_G1365 = ~new_G326;
  assign new_G1405 = new_G401;
  assign new_G285 = ~new_G279;
  assign new_G347 = ~new_G1134 | ~new_G1143;
  assign new_G367 = ~new_G366;
  assign new_G415 = ~new_G413 | ~new_G414;
  assign new_G1393 = ~new_G1389;
  assign new_G556 = ~new_G1501 | ~new_G1504;
  assign new_G1505 = ~new_G1501;
  assign new_G559 = ~new_G1493 | ~new_G1496;
  assign new_G1497 = ~new_G1493;
  assign new_G1693 = ~new_G1689;
  assign new_G1133 = ~new_G1122 | ~new_G1131;
  assign new_G1477 = new_G445;
  assign new_G1485 = new_G445;
  assign new_G1809 = ~new_G1350 | ~new_G1351;
  assign new_G348 = ~new_G346 | ~new_G347;
  assign new_G1369 = ~new_G1365;
  assign new_G1409 = ~new_G1405;
  assign new_G557 = ~new_G1498 | ~new_G1505;
  assign new_G560 = ~new_G1490 | ~new_G1497;
  assign new_G1362 = new_G282;
  assign new_G1378 = ~new_G415;
  assign new_G1429 = new_G453;
  assign new_G1437 = new_G453;
  assign new_G1686 = new_G282;
  assign new_G1774 = ~new_G1132 | ~new_G1133;
  assign new_G1910 = new_G285 & new_G853;
  assign new_G1918 = new_G856 & new_G367;
  assign new_G544 = ~new_G1485 | ~new_G1488;
  assign new_G1489 = ~new_G1485;
  assign new_G547 = ~new_G1477 | ~new_G1480;
  assign new_G1481 = ~new_G1477;
  assign new_G558 = ~new_G556 | ~new_G557;
  assign new_G561 = ~new_G559 | ~new_G560;
  assign new_G1813 = ~new_G1809;
  assign new_G1370 = ~new_G348;
  assign new_G1368 = ~new_G1362;
  assign new_G417 = ~new_G1362 | ~new_G1369;
  assign new_G1384 = ~new_G1378;
  assign new_G424 = ~new_G1378 | ~new_G1385;
  assign new_G508 = ~new_G1437 | ~new_G1440;
  assign new_G1441 = ~new_G1437;
  assign new_G511 = ~new_G1429 | ~new_G1432;
  assign new_G1433 = ~new_G1429;
  assign new_G545 = ~new_G1482 | ~new_G1489;
  assign new_G548 = ~new_G1474 | ~new_G1481;
  assign new_G564 = ~new_G558;
  assign new_G1692 = ~new_G1686;
  assign new_G1024 = ~new_G1686 | ~new_G1693;
  assign new_G1780 = ~new_G1774;
  assign new_G1148 = ~new_G1774 | ~new_G1781;
  assign new_G1916 = ~new_G1910;
  assign new_G1924 = ~new_G1918;
  assign new_G416 = ~new_G1365 | ~new_G1368;
  assign new_G1376 = ~new_G1370;
  assign new_G421 = ~new_G1370 | ~new_G1377;
  assign new_G423 = ~new_G1381 | ~new_G1384;
  assign new_G509 = ~new_G1434 | ~new_G1441;
  assign new_G512 = ~new_G1426 | ~new_G1433;
  assign new_G546 = ~new_G544 | ~new_G545;
  assign new_G549 = ~new_G547 | ~new_G548;
  assign new_G719 = ~new_G561;
  assign new_G722 = new_G561;
  assign new_G1023 = ~new_G1689 | ~new_G1692;
  assign new_G1147 = ~new_G1777 | ~new_G1780;
  assign new_G418 = ~new_G416 | ~new_G417;
  assign new_G420 = ~new_G1373 | ~new_G1376;
  assign new_G425 = ~new_G423 | ~new_G424;
  assign new_G510 = ~new_G508 | ~new_G509;
  assign new_G513 = ~new_G511 | ~new_G512;
  assign new_G552 = ~new_G546;
  assign new_G1025 = ~new_G1023 | ~new_G1024;
  assign new_G1149 = ~new_G1147 | ~new_G1148;
  assign new_G419 = ~new_G418;
  assign new_G422 = ~new_G420 | ~new_G421;
  assign new_G441 = ~new_G425 | ~new_G918;
  assign new_G516 = ~new_G510;
  assign new_G725 = ~new_G549;
  assign new_G728 = new_G549;
  assign new_G1029 = ~new_G1025;
  assign new_G1153 = ~new_G1149;
  assign new_G433 = ~new_G419 | ~new_G918;
  assign new_G437 = ~new_G422 | ~new_G918;
  assign new_G663 = ~new_G513;
  assign new_G666 = new_G513;
  assign new_G731 = new_G719 & new_G725;
  assign new_G746 = new_G722 & new_G725;
  assign new_G756 = new_G719 & new_G728;
  assign new_G770 = new_G722 & new_G728;
  assign new_G1461 = new_G441;
  assign new_G1469 = new_G441;
  assign new_G1413 = new_G433;
  assign new_G1421 = new_G433;
  assign new_G1445 = new_G437;
  assign new_G1453 = new_G437;
  assign new_G532 = ~new_G1469 | ~new_G1472;
  assign new_G1473 = ~new_G1469;
  assign new_G535 = ~new_G1461 | ~new_G1464;
  assign new_G1465 = ~new_G1461;
  assign new_G495 = ~new_G1421 | ~new_G1424;
  assign new_G1425 = ~new_G1421;
  assign new_G498 = ~new_G1413 | ~new_G1416;
  assign new_G1417 = ~new_G1413;
  assign new_G520 = ~new_G1453 | ~new_G1456;
  assign new_G1457 = ~new_G1453;
  assign new_G523 = ~new_G1445 | ~new_G1448;
  assign new_G1449 = ~new_G1445;
  assign new_G533 = ~new_G1466 | ~new_G1473;
  assign new_G536 = ~new_G1458 | ~new_G1465;
  assign new_G496 = ~new_G1418 | ~new_G1425;
  assign new_G499 = ~new_G1410 | ~new_G1417;
  assign new_G521 = ~new_G1450 | ~new_G1457;
  assign new_G524 = ~new_G1442 | ~new_G1449;
  assign new_G534 = ~new_G532 | ~new_G533;
  assign new_G537 = ~new_G535 | ~new_G536;
  assign new_G497 = ~new_G495 | ~new_G496;
  assign new_G500 = ~new_G498 | ~new_G499;
  assign new_G522 = ~new_G520 | ~new_G521;
  assign new_G525 = ~new_G523 | ~new_G524;
  assign new_G540 = ~new_G534;
  assign new_G503 = ~new_G497;
  assign new_G528 = ~new_G522;
  assign new_G669 = ~new_G537;
  assign new_G672 = new_G537;
  assign new_G569 = ~new_G500;
  assign new_G588 = new_G566 & new_G500;
  assign new_G618 = ~new_G525;
  assign new_G639 = new_G615 & new_G525;
  assign new_G867 = ~new_G487 | ~new_G503 | ~new_G528 | ~new_G482 | ~new_G540 | ~new_G552 | ~new_G516 | ~new_G564;
  assign new_G588a = new_G588;
  assign new_G588b = new_G588;
  assign new_G639a = new_G639;
  assign new_G639b = new_G639;
  assign new_G675 = new_G663 & new_G669;
  assign new_G688 = new_G666 & new_G669;
  assign new_G696 = new_G663 & new_G672;
  assign new_G710 = new_G666 & new_G672;
  assign new_G73 = new_G932 & new_G932 & new_G949 & new_G867;
  assign new_G572 = new_G565 & new_G569;
  assign new_G573 = new_G566 & new_G569;
  assign new_G621 = new_G614 & new_G618;
  assign new_G622 = new_G615 & new_G618;
  assign new_G776 = ~new_G958 | ~new_G731 | ~new_G696 | ~new_G588a | ~new_G639a;
  assign new_G780 = ~new_G958 | ~new_G756 | ~new_G675 | ~new_G588a | ~new_G639a;
  assign new_G784 = ~new_G958 | ~new_G746 | ~new_G675 | ~new_G588a | ~new_G639a;
  assign new_G788 = ~new_G958 | ~new_G731 | ~new_G688 | ~new_G588a | ~new_G639a;
  assign new_G812 = ~new_G969 | ~new_G746 | ~new_G710 | ~new_G588b | ~new_G639a;
  assign new_G832 = ~new_G969 | ~new_G770 | ~new_G696 | ~new_G588b | ~new_G639b;
  assign new_G836 = ~new_G969 | ~new_G756 | ~new_G710 | ~new_G588b | ~new_G639b;
  assign new_G1509 = new_G958 & new_G731 & new_G696 & new_G588a & new_G639a;
  assign new_G1517 = new_G958 & new_G756 & new_G675 & new_G588a & new_G639a;
  assign new_G1525 = new_G958 & new_G746 & new_G675 & new_G588a & new_G639a;
  assign new_G1533 = new_G958 & new_G731 & new_G688 & new_G588a & new_G639a;
  assign new_G1581 = new_G969 & new_G746 & new_G710 & new_G588b & new_G639a;
  assign new_G1621 = new_G969 & new_G770 & new_G696 & new_G588b & new_G639b;
  assign new_G1629 = new_G969 & new_G756 & new_G710 & new_G588b & new_G639b;
  assign new_G792 = ~new_G958 | ~new_G756 | ~new_G696 | ~new_G588a | ~new_G622;
  assign new_G796 = ~new_G958 | ~new_G746 | ~new_G696 | ~new_G588b | ~new_G622;
  assign new_G800 = ~new_G958 | ~new_G731 | ~new_G710 | ~new_G588b | ~new_G622;
  assign new_G804 = ~new_G958 | ~new_G770 | ~new_G675 | ~new_G588b | ~new_G622;
  assign new_G808 = ~new_G969 | ~new_G756 | ~new_G688 | ~new_G588b | ~new_G622;
  assign new_G816 = ~new_G969 | ~new_G756 | ~new_G696 | ~new_G573 | ~new_G639b;
  assign new_G820 = ~new_G969 | ~new_G746 | ~new_G696 | ~new_G573 | ~new_G639b;
  assign new_G824 = ~new_G969 | ~new_G731 | ~new_G710 | ~new_G573 | ~new_G639b;
  assign new_G828 = ~new_G969 | ~new_G756 | ~new_G688 | ~new_G573 | ~new_G639b;
  assign new_G871 = ~new_G979 | ~new_G731 | ~new_G675 | ~new_G588b | ~new_G622;
  assign new_G873 = ~new_G979 | ~new_G731 | ~new_G675 | ~new_G573 | ~new_G639b;
  assign new_G875 = ~new_G979 | ~new_G731 | ~new_G696 | ~new_G573 | ~new_G622;
  assign new_G877 = ~new_G979 | ~new_G756 | ~new_G675 | ~new_G573 | ~new_G622;
  assign new_G879 = ~new_G979 | ~new_G746 | ~new_G675 | ~new_G573 | ~new_G622;
  assign new_G881 = ~new_G979 | ~new_G731 | ~new_G688 | ~new_G573 | ~new_G622;
  assign new_G883 = ~new_G979 | ~new_G731 | ~new_G675 | ~new_G573 | ~new_G621;
  assign new_G885 = ~new_G979 | ~new_G731 | ~new_G675 | ~new_G572 | ~new_G622;
  assign new_G1541 = new_G958 & new_G756 & new_G696 & new_G588a & new_G622;
  assign new_G1549 = new_G958 & new_G746 & new_G696 & new_G588b & new_G622;
  assign new_G1557 = new_G958 & new_G731 & new_G710 & new_G588b & new_G622;
  assign new_G1565 = new_G958 & new_G770 & new_G675 & new_G588b & new_G622;
  assign new_G1573 = new_G969 & new_G756 & new_G688 & new_G588b & new_G622;
  assign new_G1589 = new_G969 & new_G756 & new_G696 & new_G573 & new_G639b;
  assign new_G1597 = new_G969 & new_G746 & new_G696 & new_G573 & new_G639b;
  assign new_G1605 = new_G969 & new_G731 & new_G710 & new_G573 & new_G639b;
  assign new_G1613 = new_G969 & new_G756 & new_G688 & new_G573 & new_G639b;
  assign new_G1 = ~new_G1509 | ~new_G1512;
  assign new_G1513 = ~new_G1509;
  assign new_G4 = ~new_G1517 | ~new_G1520;
  assign new_G1521 = ~new_G1517;
  assign new_G7 = ~new_G1525 | ~new_G1528;
  assign new_G1529 = ~new_G1525;
  assign new_G10 = ~new_G1533 | ~new_G1536;
  assign new_G1537 = ~new_G1533;
  assign new_G28 = ~new_G1581 | ~new_G1584;
  assign new_G1585 = ~new_G1581;
  assign new_G43 = ~new_G1621 | ~new_G1624;
  assign new_G1625 = ~new_G1621;
  assign new_G46 = ~new_G1629 | ~new_G1632;
  assign new_G1633 = ~new_G1629;
  assign new_G886 = new_G885 & new_G883 & new_G881 & new_G879 & new_G877 & new_G875 & new_G871 & new_G873;
  assign new_G2 = ~new_G1506 | ~new_G1513;
  assign new_G5 = ~new_G1514 | ~new_G1521;
  assign new_G8 = ~new_G1522 | ~new_G1529;
  assign new_G11 = ~new_G1530 | ~new_G1537;
  assign new_G13 = ~new_G1541 | ~new_G1544;
  assign new_G1545 = ~new_G1541;
  assign new_G16 = ~new_G1549 | ~new_G1552;
  assign new_G1553 = ~new_G1549;
  assign new_G19 = ~new_G1557 | ~new_G1560;
  assign new_G1561 = ~new_G1557;
  assign new_G22 = ~new_G1565 | ~new_G1568;
  assign new_G1569 = ~new_G1565;
  assign new_G25 = ~new_G1573 | ~new_G1576;
  assign new_G1577 = ~new_G1573;
  assign new_G29 = ~new_G1578 | ~new_G1585;
  assign new_G31 = ~new_G1589 | ~new_G1592;
  assign new_G1593 = ~new_G1589;
  assign new_G34 = ~new_G1597 | ~new_G1600;
  assign new_G1601 = ~new_G1597;
  assign new_G37 = ~new_G1605 | ~new_G1608;
  assign new_G1609 = ~new_G1605;
  assign new_G40 = ~new_G1613 | ~new_G1616;
  assign new_G1617 = ~new_G1613;
  assign new_G44 = ~new_G1618 | ~new_G1625;
  assign new_G47 = ~new_G1626 | ~new_G1633;
  assign new_G857 = ~new_G804 | ~new_G800 | ~new_G796 | ~new_G792 | ~new_G788 | ~new_G784 | ~new_G776 | ~new_G780;
  assign new_G860 = ~new_G836 | ~new_G832 | ~new_G828 | ~new_G824 | ~new_G820 | ~new_G816 | ~new_G808 | ~new_G812;
  assign new_G863 = new_G804 & new_G800 & new_G796 & new_G792 & new_G788 & new_G784 & new_G776 & new_G780;
  assign new_G865 = new_G836 & new_G832 & new_G828 & new_G824 & new_G820 & new_G816 & new_G808 & new_G812;
  assign G3 = ~new_G1 | ~new_G2;
  assign G6 = ~new_G4 | ~new_G5;
  assign G9 = ~new_G7 | ~new_G8;
  assign G12 = ~new_G10 | ~new_G11;
  assign new_G14 = ~new_G1538 | ~new_G1545;
  assign new_G17 = ~new_G1546 | ~new_G1553;
  assign new_G20 = ~new_G1554 | ~new_G1561;
  assign new_G23 = ~new_G1562 | ~new_G1569;
  assign new_G26 = ~new_G1570 | ~new_G1577;
  assign G30 = ~new_G28 | ~new_G29;
  assign new_G32 = ~new_G1586 | ~new_G1593;
  assign new_G35 = ~new_G1594 | ~new_G1601;
  assign new_G38 = ~new_G1602 | ~new_G1609;
  assign new_G41 = ~new_G1610 | ~new_G1617;
  assign G45 = ~new_G43 | ~new_G44;
  assign G48 = ~new_G46 | ~new_G47;
  assign new_G1913 = new_G857 & new_G859;
  assign new_G1921 = new_G860 & new_G862;
  assign G15 = ~new_G13 | ~new_G14;
  assign G18 = ~new_G16 | ~new_G17;
  assign G21 = ~new_G19 | ~new_G20;
  assign G24 = ~new_G22 | ~new_G23;
  assign G27 = ~new_G25 | ~new_G26;
  assign G33 = ~new_G31 | ~new_G32;
  assign G36 = ~new_G34 | ~new_G35;
  assign G39 = ~new_G37 | ~new_G38;
  assign G42 = ~new_G40 | ~new_G41;
  assign new_G887 = new_G886 & new_G863 & new_G865;
  assign new_G462 = ~new_G863 | ~new_G865;
  assign new_G74 = new_G887 & G952 & new_G949 & new_G867;
  assign new_G1637 = ~new_G1913 | ~new_G1916;
  assign new_G1917 = ~new_G1913;
  assign new_G1647 = ~new_G1921 | ~new_G1924;
  assign new_G1925 = ~new_G1921;
  assign G75 = ~new_G73 & ~new_G74;
  assign new_G1020 = new_G462 & new_G457 & new_G911;
  assign new_G1144 = new_G462 & G469 & new_G911;
  assign new_G1386 = new_G462 & G475 & new_G911;
  assign new_G1394 = new_G462 & G478 & new_G911;
  assign new_G1402 = new_G462 & new_G459 & new_G911;
  assign new_G1638 = ~new_G1910 | ~new_G1917;
  assign new_G1648 = ~new_G1918 | ~new_G1925;
  assign new_G1806 = new_G462 & G472 & new_G911;
  assign new_G1639 = ~new_G1637 | ~new_G1638;
  assign new_G1649 = ~new_G1647 | ~new_G1648;
  assign new_G287 = ~new_G1020 | ~new_G1029;
  assign new_G350 = ~new_G1144 | ~new_G1153;
  assign new_G427 = ~new_G1386 | ~new_G1393;
  assign new_G429 = ~new_G1394 | ~new_G1401;
  assign new_G431 = ~new_G1402 | ~new_G1409;
  assign new_G1028 = ~new_G1020;
  assign new_G1152 = ~new_G1144;
  assign new_G1392 = ~new_G1386;
  assign new_G1400 = ~new_G1394;
  assign new_G1408 = ~new_G1402;
  assign new_G1812 = ~new_G1806;
  assign new_G1216 = ~new_G1806 | ~new_G1813;
  assign new_G286 = ~new_G1025 | ~new_G1028;
  assign new_G349 = ~new_G1149 | ~new_G1152;
  assign new_G426 = ~new_G1389 | ~new_G1392;
  assign new_G428 = ~new_G1397 | ~new_G1400;
  assign new_G430 = ~new_G1405 | ~new_G1408;
  assign new_G67 = ~new_G1639 | ~new_G1642;
  assign new_G1643 = ~new_G1639;
  assign new_G70 = ~new_G1649 | ~new_G1652;
  assign new_G1653 = ~new_G1649;
  assign new_G1215 = ~new_G1809 | ~new_G1812;
  assign new_G49 = ~new_G286 | ~new_G287;
  assign new_G53 = ~new_G349 | ~new_G350;
  assign new_G59 = ~new_G426 | ~new_G427;
  assign new_G61 = ~new_G428 | ~new_G429;
  assign new_G65 = ~new_G430 | ~new_G431;
  assign new_G68 = ~new_G1634 | ~new_G1643;
  assign new_G71 = ~new_G1644 | ~new_G1653;
  assign new_G1217 = ~new_G1215 | ~new_G1216;
  assign G51 = new_G49 & new_G50;
  assign G54 = new_G52 & new_G53;
  assign G60 = new_G58 & new_G59;
  assign G63 = new_G61 & new_G62;
  assign G66 = new_G64 & new_G65;
  assign G69 = ~new_G67 | ~new_G68;
  assign G72 = ~new_G70 | ~new_G71;
  assign new_G375 = ~new_G1217 | ~new_G1220;
  assign new_G1221 = ~new_G1217;
  assign new_G376 = ~new_G1212 | ~new_G1221;
  assign new_G55 = ~new_G375 | ~new_G376;
  assign G57 = new_G55 & new_G56;
endmodule
